module IssueUnitCollapsing_2(
  input         clock,
  input         reset,
  output        io_dis_uops_0_ready,
  input         io_dis_uops_0_valid,
  input         io_dis_uops_0_bits_switch,
  input         io_dis_uops_0_bits_switch_off,
  input         io_dis_uops_0_bits_is_unicore,
  input  [2:0]  io_dis_uops_0_bits_shift,
  input  [1:0]  io_dis_uops_0_bits_lrs3_rtype,
  input         io_dis_uops_0_bits_rflag,
  input         io_dis_uops_0_bits_wflag,
  input  [3:0]  io_dis_uops_0_bits_prflag,
  input  [3:0]  io_dis_uops_0_bits_pwflag,
  input         io_dis_uops_0_bits_pflag_busy,
  input  [3:0]  io_dis_uops_0_bits_stale_pflag,
  input  [3:0]  io_dis_uops_0_bits_op1_sel,
  input  [3:0]  io_dis_uops_0_bits_op2_sel,
  input  [5:0]  io_dis_uops_0_bits_split_num,
  input  [5:0]  io_dis_uops_0_bits_self_index,
  input  [5:0]  io_dis_uops_0_bits_rob_inst_idx,
  input  [5:0]  io_dis_uops_0_bits_address_num,
  input  [6:0]  io_dis_uops_0_bits_uopc,
  input  [31:0] io_dis_uops_0_bits_inst,
  input  [31:0] io_dis_uops_0_bits_debug_inst,
  input         io_dis_uops_0_bits_is_rvc,
  input  [39:0] io_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_dis_uops_0_bits_iq_type,
  input  [9:0]  io_dis_uops_0_bits_fu_code,
  input  [3:0]  io_dis_uops_0_bits_ctrl_br_type,
  input  [1:0]  io_dis_uops_0_bits_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_0_bits_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_0_bits_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_0_bits_ctrl_op_fcn,
  input         io_dis_uops_0_bits_ctrl_fcn_dw,
  input  [2:0]  io_dis_uops_0_bits_ctrl_csr_cmd,
  input         io_dis_uops_0_bits_ctrl_is_load,
  input         io_dis_uops_0_bits_ctrl_is_sta,
  input         io_dis_uops_0_bits_ctrl_is_std,
  input  [1:0]  io_dis_uops_0_bits_ctrl_op3_sel,
  input  [1:0]  io_dis_uops_0_bits_iw_state,
  input         io_dis_uops_0_bits_iw_p1_poisoned,
  input         io_dis_uops_0_bits_iw_p2_poisoned,
  input         io_dis_uops_0_bits_is_br,
  input         io_dis_uops_0_bits_is_jalr,
  input         io_dis_uops_0_bits_is_jal,
  input         io_dis_uops_0_bits_is_sfb,
  input  [11:0] io_dis_uops_0_bits_br_mask,
  input  [3:0]  io_dis_uops_0_bits_br_tag,
  input  [4:0]  io_dis_uops_0_bits_ftq_idx,
  input         io_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_dis_uops_0_bits_pc_lob,
  input         io_dis_uops_0_bits_taken,
  input  [19:0] io_dis_uops_0_bits_imm_packed,
  input  [11:0] io_dis_uops_0_bits_csr_addr,
  input  [5:0]  io_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_dis_uops_0_bits_ldq_idx,
  input  [4:0]  io_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_dis_uops_0_bits_pdst,
  input  [6:0]  io_dis_uops_0_bits_prs1,
  input  [6:0]  io_dis_uops_0_bits_prs2,
  input  [6:0]  io_dis_uops_0_bits_prs3,
  input  [4:0]  io_dis_uops_0_bits_ppred,
  input         io_dis_uops_0_bits_prs1_busy,
  input         io_dis_uops_0_bits_prs2_busy,
  input         io_dis_uops_0_bits_prs3_busy,
  input         io_dis_uops_0_bits_ppred_busy,
  input  [6:0]  io_dis_uops_0_bits_stale_pdst,
  input         io_dis_uops_0_bits_exception,
  input  [63:0] io_dis_uops_0_bits_exc_cause,
  input         io_dis_uops_0_bits_bypassable,
  input  [4:0]  io_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_dis_uops_0_bits_mem_size,
  input         io_dis_uops_0_bits_mem_signed,
  input         io_dis_uops_0_bits_is_fence,
  input         io_dis_uops_0_bits_is_fencei,
  input         io_dis_uops_0_bits_is_amo,
  input         io_dis_uops_0_bits_uses_ldq,
  input         io_dis_uops_0_bits_uses_stq,
  input         io_dis_uops_0_bits_is_sys_pc2epc,
  input         io_dis_uops_0_bits_is_unique,
  input         io_dis_uops_0_bits_flush_on_commit,
  input         io_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_0_bits_ldst,
  input  [5:0]  io_dis_uops_0_bits_lrs1,
  input  [5:0]  io_dis_uops_0_bits_lrs2,
  input  [5:0]  io_dis_uops_0_bits_lrs3,
  input         io_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_dis_uops_0_bits_dst_rtype,
  input  [1:0]  io_dis_uops_0_bits_lrs1_rtype,
  input  [1:0]  io_dis_uops_0_bits_lrs2_rtype,
  input         io_dis_uops_0_bits_frs3_en,
  input         io_dis_uops_0_bits_fp_val,
  input         io_dis_uops_0_bits_fp_single,
  input         io_dis_uops_0_bits_xcpt_pf_if,
  input         io_dis_uops_0_bits_xcpt_ae_if,
  input         io_dis_uops_0_bits_xcpt_ma_if,
  input         io_dis_uops_0_bits_bp_debug_if,
  input         io_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_0_bits_debug_fsrc,
  input  [1:0]  io_dis_uops_0_bits_debug_tsrc,
  output        io_dis_uops_1_ready,
  input         io_dis_uops_1_valid,
  input         io_dis_uops_1_bits_switch,
  input         io_dis_uops_1_bits_switch_off,
  input         io_dis_uops_1_bits_is_unicore,
  input  [2:0]  io_dis_uops_1_bits_shift,
  input  [1:0]  io_dis_uops_1_bits_lrs3_rtype,
  input         io_dis_uops_1_bits_rflag,
  input         io_dis_uops_1_bits_wflag,
  input  [3:0]  io_dis_uops_1_bits_prflag,
  input  [3:0]  io_dis_uops_1_bits_pwflag,
  input         io_dis_uops_1_bits_pflag_busy,
  input  [3:0]  io_dis_uops_1_bits_stale_pflag,
  input  [3:0]  io_dis_uops_1_bits_op1_sel,
  input  [3:0]  io_dis_uops_1_bits_op2_sel,
  input  [5:0]  io_dis_uops_1_bits_split_num,
  input  [5:0]  io_dis_uops_1_bits_self_index,
  input  [5:0]  io_dis_uops_1_bits_rob_inst_idx,
  input  [5:0]  io_dis_uops_1_bits_address_num,
  input  [6:0]  io_dis_uops_1_bits_uopc,
  input  [31:0] io_dis_uops_1_bits_inst,
  input  [31:0] io_dis_uops_1_bits_debug_inst,
  input         io_dis_uops_1_bits_is_rvc,
  input  [39:0] io_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_dis_uops_1_bits_iq_type,
  input  [9:0]  io_dis_uops_1_bits_fu_code,
  input  [3:0]  io_dis_uops_1_bits_ctrl_br_type,
  input  [1:0]  io_dis_uops_1_bits_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_1_bits_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_1_bits_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_1_bits_ctrl_op_fcn,
  input         io_dis_uops_1_bits_ctrl_fcn_dw,
  input  [2:0]  io_dis_uops_1_bits_ctrl_csr_cmd,
  input         io_dis_uops_1_bits_ctrl_is_load,
  input         io_dis_uops_1_bits_ctrl_is_sta,
  input         io_dis_uops_1_bits_ctrl_is_std,
  input  [1:0]  io_dis_uops_1_bits_ctrl_op3_sel,
  input  [1:0]  io_dis_uops_1_bits_iw_state,
  input         io_dis_uops_1_bits_iw_p1_poisoned,
  input         io_dis_uops_1_bits_iw_p2_poisoned,
  input         io_dis_uops_1_bits_is_br,
  input         io_dis_uops_1_bits_is_jalr,
  input         io_dis_uops_1_bits_is_jal,
  input         io_dis_uops_1_bits_is_sfb,
  input  [11:0] io_dis_uops_1_bits_br_mask,
  input  [3:0]  io_dis_uops_1_bits_br_tag,
  input  [4:0]  io_dis_uops_1_bits_ftq_idx,
  input         io_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_dis_uops_1_bits_pc_lob,
  input         io_dis_uops_1_bits_taken,
  input  [19:0] io_dis_uops_1_bits_imm_packed,
  input  [11:0] io_dis_uops_1_bits_csr_addr,
  input  [5:0]  io_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_dis_uops_1_bits_ldq_idx,
  input  [4:0]  io_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_dis_uops_1_bits_pdst,
  input  [6:0]  io_dis_uops_1_bits_prs1,
  input  [6:0]  io_dis_uops_1_bits_prs2,
  input  [6:0]  io_dis_uops_1_bits_prs3,
  input  [4:0]  io_dis_uops_1_bits_ppred,
  input         io_dis_uops_1_bits_prs1_busy,
  input         io_dis_uops_1_bits_prs2_busy,
  input         io_dis_uops_1_bits_prs3_busy,
  input         io_dis_uops_1_bits_ppred_busy,
  input  [6:0]  io_dis_uops_1_bits_stale_pdst,
  input         io_dis_uops_1_bits_exception,
  input  [63:0] io_dis_uops_1_bits_exc_cause,
  input         io_dis_uops_1_bits_bypassable,
  input  [4:0]  io_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_dis_uops_1_bits_mem_size,
  input         io_dis_uops_1_bits_mem_signed,
  input         io_dis_uops_1_bits_is_fence,
  input         io_dis_uops_1_bits_is_fencei,
  input         io_dis_uops_1_bits_is_amo,
  input         io_dis_uops_1_bits_uses_ldq,
  input         io_dis_uops_1_bits_uses_stq,
  input         io_dis_uops_1_bits_is_sys_pc2epc,
  input         io_dis_uops_1_bits_is_unique,
  input         io_dis_uops_1_bits_flush_on_commit,
  input         io_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_1_bits_ldst,
  input  [5:0]  io_dis_uops_1_bits_lrs1,
  input  [5:0]  io_dis_uops_1_bits_lrs2,
  input  [5:0]  io_dis_uops_1_bits_lrs3,
  input         io_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_dis_uops_1_bits_dst_rtype,
  input  [1:0]  io_dis_uops_1_bits_lrs1_rtype,
  input  [1:0]  io_dis_uops_1_bits_lrs2_rtype,
  input         io_dis_uops_1_bits_frs3_en,
  input         io_dis_uops_1_bits_fp_val,
  input         io_dis_uops_1_bits_fp_single,
  input         io_dis_uops_1_bits_xcpt_pf_if,
  input         io_dis_uops_1_bits_xcpt_ae_if,
  input         io_dis_uops_1_bits_xcpt_ma_if,
  input         io_dis_uops_1_bits_bp_debug_if,
  input         io_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_1_bits_debug_fsrc,
  input  [1:0]  io_dis_uops_1_bits_debug_tsrc,
  output        io_iss_valids_0,
  output        io_iss_valids_1,
  output        io_iss_uops_0_switch,
  output        io_iss_uops_0_switch_off,
  output        io_iss_uops_0_is_unicore,
  output [2:0]  io_iss_uops_0_shift,
  output [1:0]  io_iss_uops_0_lrs3_rtype,
  output        io_iss_uops_0_rflag,
  output        io_iss_uops_0_wflag,
  output [3:0]  io_iss_uops_0_prflag,
  output [3:0]  io_iss_uops_0_pwflag,
  output        io_iss_uops_0_pflag_busy,
  output [3:0]  io_iss_uops_0_stale_pflag,
  output [3:0]  io_iss_uops_0_op1_sel,
  output [3:0]  io_iss_uops_0_op2_sel,
  output [5:0]  io_iss_uops_0_split_num,
  output [5:0]  io_iss_uops_0_self_index,
  output [5:0]  io_iss_uops_0_rob_inst_idx,
  output [5:0]  io_iss_uops_0_address_num,
  output [6:0]  io_iss_uops_0_uopc,
  output [31:0] io_iss_uops_0_inst,
  output [31:0] io_iss_uops_0_debug_inst,
  output        io_iss_uops_0_is_rvc,
  output [39:0] io_iss_uops_0_debug_pc,
  output [2:0]  io_iss_uops_0_iq_type,
  output [9:0]  io_iss_uops_0_fu_code,
  output [3:0]  io_iss_uops_0_ctrl_br_type,
  output [1:0]  io_iss_uops_0_ctrl_op1_sel,
  output [2:0]  io_iss_uops_0_ctrl_op2_sel,
  output [2:0]  io_iss_uops_0_ctrl_imm_sel,
  output [3:0]  io_iss_uops_0_ctrl_op_fcn,
  output        io_iss_uops_0_ctrl_fcn_dw,
  output [2:0]  io_iss_uops_0_ctrl_csr_cmd,
  output        io_iss_uops_0_ctrl_is_load,
  output        io_iss_uops_0_ctrl_is_sta,
  output        io_iss_uops_0_ctrl_is_std,
  output [1:0]  io_iss_uops_0_ctrl_op3_sel,
  output [1:0]  io_iss_uops_0_iw_state,
  output        io_iss_uops_0_iw_p1_poisoned,
  output        io_iss_uops_0_iw_p2_poisoned,
  output        io_iss_uops_0_is_br,
  output        io_iss_uops_0_is_jalr,
  output        io_iss_uops_0_is_jal,
  output        io_iss_uops_0_is_sfb,
  output [11:0] io_iss_uops_0_br_mask,
  output [3:0]  io_iss_uops_0_br_tag,
  output [4:0]  io_iss_uops_0_ftq_idx,
  output        io_iss_uops_0_edge_inst,
  output [5:0]  io_iss_uops_0_pc_lob,
  output        io_iss_uops_0_taken,
  output [19:0] io_iss_uops_0_imm_packed,
  output [11:0] io_iss_uops_0_csr_addr,
  output [5:0]  io_iss_uops_0_rob_idx,
  output [4:0]  io_iss_uops_0_ldq_idx,
  output [4:0]  io_iss_uops_0_stq_idx,
  output [1:0]  io_iss_uops_0_rxq_idx,
  output [6:0]  io_iss_uops_0_pdst,
  output [6:0]  io_iss_uops_0_prs1,
  output [6:0]  io_iss_uops_0_prs2,
  output [6:0]  io_iss_uops_0_prs3,
  output [4:0]  io_iss_uops_0_ppred,
  output        io_iss_uops_0_prs1_busy,
  output        io_iss_uops_0_prs2_busy,
  output        io_iss_uops_0_prs3_busy,
  output        io_iss_uops_0_ppred_busy,
  output [6:0]  io_iss_uops_0_stale_pdst,
  output        io_iss_uops_0_exception,
  output [63:0] io_iss_uops_0_exc_cause,
  output        io_iss_uops_0_bypassable,
  output [4:0]  io_iss_uops_0_mem_cmd,
  output [1:0]  io_iss_uops_0_mem_size,
  output        io_iss_uops_0_mem_signed,
  output        io_iss_uops_0_is_fence,
  output        io_iss_uops_0_is_fencei,
  output        io_iss_uops_0_is_amo,
  output        io_iss_uops_0_uses_ldq,
  output        io_iss_uops_0_uses_stq,
  output        io_iss_uops_0_is_sys_pc2epc,
  output        io_iss_uops_0_is_unique,
  output        io_iss_uops_0_flush_on_commit,
  output        io_iss_uops_0_ldst_is_rs1,
  output [5:0]  io_iss_uops_0_ldst,
  output [5:0]  io_iss_uops_0_lrs1,
  output [5:0]  io_iss_uops_0_lrs2,
  output [5:0]  io_iss_uops_0_lrs3,
  output        io_iss_uops_0_ldst_val,
  output [1:0]  io_iss_uops_0_dst_rtype,
  output [1:0]  io_iss_uops_0_lrs1_rtype,
  output [1:0]  io_iss_uops_0_lrs2_rtype,
  output        io_iss_uops_0_frs3_en,
  output        io_iss_uops_0_fp_val,
  output        io_iss_uops_0_fp_single,
  output        io_iss_uops_0_xcpt_pf_if,
  output        io_iss_uops_0_xcpt_ae_if,
  output        io_iss_uops_0_xcpt_ma_if,
  output        io_iss_uops_0_bp_debug_if,
  output        io_iss_uops_0_bp_xcpt_if,
  output [1:0]  io_iss_uops_0_debug_fsrc,
  output [1:0]  io_iss_uops_0_debug_tsrc,
  output        io_iss_uops_1_switch,
  output        io_iss_uops_1_switch_off,
  output        io_iss_uops_1_is_unicore,
  output [2:0]  io_iss_uops_1_shift,
  output [1:0]  io_iss_uops_1_lrs3_rtype,
  output        io_iss_uops_1_rflag,
  output        io_iss_uops_1_wflag,
  output [3:0]  io_iss_uops_1_prflag,
  output [3:0]  io_iss_uops_1_pwflag,
  output        io_iss_uops_1_pflag_busy,
  output [3:0]  io_iss_uops_1_stale_pflag,
  output [3:0]  io_iss_uops_1_op1_sel,
  output [3:0]  io_iss_uops_1_op2_sel,
  output [5:0]  io_iss_uops_1_split_num,
  output [5:0]  io_iss_uops_1_self_index,
  output [5:0]  io_iss_uops_1_rob_inst_idx,
  output [5:0]  io_iss_uops_1_address_num,
  output [6:0]  io_iss_uops_1_uopc,
  output [31:0] io_iss_uops_1_inst,
  output [31:0] io_iss_uops_1_debug_inst,
  output        io_iss_uops_1_is_rvc,
  output [39:0] io_iss_uops_1_debug_pc,
  output [2:0]  io_iss_uops_1_iq_type,
  output [9:0]  io_iss_uops_1_fu_code,
  output [3:0]  io_iss_uops_1_ctrl_br_type,
  output [1:0]  io_iss_uops_1_ctrl_op1_sel,
  output [2:0]  io_iss_uops_1_ctrl_op2_sel,
  output [2:0]  io_iss_uops_1_ctrl_imm_sel,
  output [3:0]  io_iss_uops_1_ctrl_op_fcn,
  output        io_iss_uops_1_ctrl_fcn_dw,
  output [2:0]  io_iss_uops_1_ctrl_csr_cmd,
  output        io_iss_uops_1_ctrl_is_load,
  output        io_iss_uops_1_ctrl_is_sta,
  output        io_iss_uops_1_ctrl_is_std,
  output [1:0]  io_iss_uops_1_ctrl_op3_sel,
  output [1:0]  io_iss_uops_1_iw_state,
  output        io_iss_uops_1_iw_p1_poisoned,
  output        io_iss_uops_1_iw_p2_poisoned,
  output        io_iss_uops_1_is_br,
  output        io_iss_uops_1_is_jalr,
  output        io_iss_uops_1_is_jal,
  output        io_iss_uops_1_is_sfb,
  output [11:0] io_iss_uops_1_br_mask,
  output [3:0]  io_iss_uops_1_br_tag,
  output [4:0]  io_iss_uops_1_ftq_idx,
  output        io_iss_uops_1_edge_inst,
  output [5:0]  io_iss_uops_1_pc_lob,
  output        io_iss_uops_1_taken,
  output [19:0] io_iss_uops_1_imm_packed,
  output [11:0] io_iss_uops_1_csr_addr,
  output [5:0]  io_iss_uops_1_rob_idx,
  output [4:0]  io_iss_uops_1_ldq_idx,
  output [4:0]  io_iss_uops_1_stq_idx,
  output [1:0]  io_iss_uops_1_rxq_idx,
  output [6:0]  io_iss_uops_1_pdst,
  output [6:0]  io_iss_uops_1_prs1,
  output [6:0]  io_iss_uops_1_prs2,
  output [6:0]  io_iss_uops_1_prs3,
  output [4:0]  io_iss_uops_1_ppred,
  output        io_iss_uops_1_prs1_busy,
  output        io_iss_uops_1_prs2_busy,
  output        io_iss_uops_1_prs3_busy,
  output        io_iss_uops_1_ppred_busy,
  output [6:0]  io_iss_uops_1_stale_pdst,
  output        io_iss_uops_1_exception,
  output [63:0] io_iss_uops_1_exc_cause,
  output        io_iss_uops_1_bypassable,
  output [4:0]  io_iss_uops_1_mem_cmd,
  output [1:0]  io_iss_uops_1_mem_size,
  output        io_iss_uops_1_mem_signed,
  output        io_iss_uops_1_is_fence,
  output        io_iss_uops_1_is_fencei,
  output        io_iss_uops_1_is_amo,
  output        io_iss_uops_1_uses_ldq,
  output        io_iss_uops_1_uses_stq,
  output        io_iss_uops_1_is_sys_pc2epc,
  output        io_iss_uops_1_is_unique,
  output        io_iss_uops_1_flush_on_commit,
  output        io_iss_uops_1_ldst_is_rs1,
  output [5:0]  io_iss_uops_1_ldst,
  output [5:0]  io_iss_uops_1_lrs1,
  output [5:0]  io_iss_uops_1_lrs2,
  output [5:0]  io_iss_uops_1_lrs3,
  output        io_iss_uops_1_ldst_val,
  output [1:0]  io_iss_uops_1_dst_rtype,
  output [1:0]  io_iss_uops_1_lrs1_rtype,
  output [1:0]  io_iss_uops_1_lrs2_rtype,
  output        io_iss_uops_1_frs3_en,
  output        io_iss_uops_1_fp_val,
  output        io_iss_uops_1_fp_single,
  output        io_iss_uops_1_xcpt_pf_if,
  output        io_iss_uops_1_xcpt_ae_if,
  output        io_iss_uops_1_xcpt_ma_if,
  output        io_iss_uops_1_bp_debug_if,
  output        io_iss_uops_1_bp_xcpt_if,
  output [1:0]  io_iss_uops_1_debug_fsrc,
  output [1:0]  io_iss_uops_1_debug_tsrc,
  input         io_wakeup_ports_0_valid,
  input  [6:0]  io_wakeup_ports_0_bits_pdst,
  input         io_wakeup_ports_0_bits_poisoned,
  input  [6:0]  io_wakeup_ports_0_bits_pwflag,
  input         io_wakeup_ports_0_bits_flag_valid,
  input         io_wakeup_ports_1_valid,
  input  [6:0]  io_wakeup_ports_1_bits_pdst,
  input         io_wakeup_ports_1_bits_poisoned,
  input  [6:0]  io_wakeup_ports_1_bits_pwflag,
  input         io_wakeup_ports_1_bits_flag_valid,
  input         io_wakeup_ports_2_valid,
  input  [6:0]  io_wakeup_ports_2_bits_pdst,
  input         io_wakeup_ports_2_bits_poisoned,
  input  [6:0]  io_wakeup_ports_2_bits_pwflag,
  input         io_wakeup_ports_2_bits_flag_valid,
  input         io_wakeup_ports_3_valid,
  input  [6:0]  io_wakeup_ports_3_bits_pdst,
  input         io_wakeup_ports_3_bits_poisoned,
  input  [6:0]  io_wakeup_ports_3_bits_pwflag,
  input         io_wakeup_ports_3_bits_flag_valid,
  input         io_wakeup_ports_4_valid,
  input  [6:0]  io_wakeup_ports_4_bits_pdst,
  input         io_wakeup_ports_4_bits_poisoned,
  input  [6:0]  io_wakeup_ports_4_bits_pwflag,
  input         io_wakeup_ports_4_bits_flag_valid,
  input         io_pred_wakeup_port_valid,
  input  [4:0]  io_pred_wakeup_port_bits,
  input         io_spec_ld_wakeup_0_valid,
  input  [6:0]  io_spec_ld_wakeup_0_bits,
  input  [9:0]  io_fu_types_0,
  input  [9:0]  io_fu_types_1,
  input  [11:0] io_brupdate_b1_resolve_mask,
  input  [11:0] io_brupdate_b1_mispredict_mask,
  input         io_brupdate_b2_uop_switch,
  input         io_brupdate_b2_uop_switch_off,
  input         io_brupdate_b2_uop_is_unicore,
  input  [2:0]  io_brupdate_b2_uop_shift,
  input  [1:0]  io_brupdate_b2_uop_lrs3_rtype,
  input         io_brupdate_b2_uop_rflag,
  input         io_brupdate_b2_uop_wflag,
  input  [3:0]  io_brupdate_b2_uop_prflag,
  input  [3:0]  io_brupdate_b2_uop_pwflag,
  input         io_brupdate_b2_uop_pflag_busy,
  input  [3:0]  io_brupdate_b2_uop_stale_pflag,
  input  [3:0]  io_brupdate_b2_uop_op1_sel,
  input  [3:0]  io_brupdate_b2_uop_op2_sel,
  input  [5:0]  io_brupdate_b2_uop_split_num,
  input  [5:0]  io_brupdate_b2_uop_self_index,
  input  [5:0]  io_brupdate_b2_uop_rob_inst_idx,
  input  [5:0]  io_brupdate_b2_uop_address_num,
  input  [6:0]  io_brupdate_b2_uop_uopc,
  input  [31:0] io_brupdate_b2_uop_inst,
  input  [31:0] io_brupdate_b2_uop_debug_inst,
  input         io_brupdate_b2_uop_is_rvc,
  input  [39:0] io_brupdate_b2_uop_debug_pc,
  input  [2:0]  io_brupdate_b2_uop_iq_type,
  input  [9:0]  io_brupdate_b2_uop_fu_code,
  input  [3:0]  io_brupdate_b2_uop_ctrl_br_type,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op1_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_op2_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_imm_sel,
  input  [3:0]  io_brupdate_b2_uop_ctrl_op_fcn,
  input         io_brupdate_b2_uop_ctrl_fcn_dw,
  input  [2:0]  io_brupdate_b2_uop_ctrl_csr_cmd,
  input         io_brupdate_b2_uop_ctrl_is_load,
  input         io_brupdate_b2_uop_ctrl_is_sta,
  input         io_brupdate_b2_uop_ctrl_is_std,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op3_sel,
  input  [1:0]  io_brupdate_b2_uop_iw_state,
  input         io_brupdate_b2_uop_iw_p1_poisoned,
  input         io_brupdate_b2_uop_iw_p2_poisoned,
  input         io_brupdate_b2_uop_is_br,
  input         io_brupdate_b2_uop_is_jalr,
  input         io_brupdate_b2_uop_is_jal,
  input         io_brupdate_b2_uop_is_sfb,
  input  [11:0] io_brupdate_b2_uop_br_mask,
  input  [3:0]  io_brupdate_b2_uop_br_tag,
  input  [4:0]  io_brupdate_b2_uop_ftq_idx,
  input         io_brupdate_b2_uop_edge_inst,
  input  [5:0]  io_brupdate_b2_uop_pc_lob,
  input         io_brupdate_b2_uop_taken,
  input  [19:0] io_brupdate_b2_uop_imm_packed,
  input  [11:0] io_brupdate_b2_uop_csr_addr,
  input  [5:0]  io_brupdate_b2_uop_rob_idx,
  input  [4:0]  io_brupdate_b2_uop_ldq_idx,
  input  [4:0]  io_brupdate_b2_uop_stq_idx,
  input  [1:0]  io_brupdate_b2_uop_rxq_idx,
  input  [6:0]  io_brupdate_b2_uop_pdst,
  input  [6:0]  io_brupdate_b2_uop_prs1,
  input  [6:0]  io_brupdate_b2_uop_prs2,
  input  [6:0]  io_brupdate_b2_uop_prs3,
  input  [4:0]  io_brupdate_b2_uop_ppred,
  input         io_brupdate_b2_uop_prs1_busy,
  input         io_brupdate_b2_uop_prs2_busy,
  input         io_brupdate_b2_uop_prs3_busy,
  input         io_brupdate_b2_uop_ppred_busy,
  input  [6:0]  io_brupdate_b2_uop_stale_pdst,
  input         io_brupdate_b2_uop_exception,
  input  [63:0] io_brupdate_b2_uop_exc_cause,
  input         io_brupdate_b2_uop_bypassable,
  input  [4:0]  io_brupdate_b2_uop_mem_cmd,
  input  [1:0]  io_brupdate_b2_uop_mem_size,
  input         io_brupdate_b2_uop_mem_signed,
  input         io_brupdate_b2_uop_is_fence,
  input         io_brupdate_b2_uop_is_fencei,
  input         io_brupdate_b2_uop_is_amo,
  input         io_brupdate_b2_uop_uses_ldq,
  input         io_brupdate_b2_uop_uses_stq,
  input         io_brupdate_b2_uop_is_sys_pc2epc,
  input         io_brupdate_b2_uop_is_unique,
  input         io_brupdate_b2_uop_flush_on_commit,
  input         io_brupdate_b2_uop_ldst_is_rs1,
  input  [5:0]  io_brupdate_b2_uop_ldst,
  input  [5:0]  io_brupdate_b2_uop_lrs1,
  input  [5:0]  io_brupdate_b2_uop_lrs2,
  input  [5:0]  io_brupdate_b2_uop_lrs3,
  input         io_brupdate_b2_uop_ldst_val,
  input  [1:0]  io_brupdate_b2_uop_dst_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs1_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs2_rtype,
  input         io_brupdate_b2_uop_frs3_en,
  input         io_brupdate_b2_uop_fp_val,
  input         io_brupdate_b2_uop_fp_single,
  input         io_brupdate_b2_uop_xcpt_pf_if,
  input         io_brupdate_b2_uop_xcpt_ae_if,
  input         io_brupdate_b2_uop_xcpt_ma_if,
  input         io_brupdate_b2_uop_bp_debug_if,
  input         io_brupdate_b2_uop_bp_xcpt_if,
  input  [1:0]  io_brupdate_b2_uop_debug_fsrc,
  input  [1:0]  io_brupdate_b2_uop_debug_tsrc,
  input         io_brupdate_b2_valid,
  input         io_brupdate_b2_mispredict,
  input         io_brupdate_b2_taken,
  input  [2:0]  io_brupdate_b2_cfi_type,
  input  [1:0]  io_brupdate_b2_pc_sel,
  input  [39:0] io_brupdate_b2_jalr_target,
  input  [31:0] io_brupdate_b2_target_offset,
  input         io_flush_pipeline,
  input         io_ld_miss,
  output        io_event_empty,
  input  [63:0] io_tsc_reg
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  slots_0_clock; // @[issue-unit.scala 157:73]
  wire  slots_0_reset; // @[issue-unit.scala 157:73]
  wire  slots_0_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_request; // @[issue-unit.scala 157:73]
  wire  slots_0_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_0_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_0_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_0_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_0_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_0_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_1_clock; // @[issue-unit.scala 157:73]
  wire  slots_1_reset; // @[issue-unit.scala 157:73]
  wire  slots_1_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_request; // @[issue-unit.scala 157:73]
  wire  slots_1_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_1_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_1_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_1_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_1_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_1_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_2_clock; // @[issue-unit.scala 157:73]
  wire  slots_2_reset; // @[issue-unit.scala 157:73]
  wire  slots_2_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_request; // @[issue-unit.scala 157:73]
  wire  slots_2_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_2_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_2_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_2_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_2_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_2_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_3_clock; // @[issue-unit.scala 157:73]
  wire  slots_3_reset; // @[issue-unit.scala 157:73]
  wire  slots_3_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_request; // @[issue-unit.scala 157:73]
  wire  slots_3_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_3_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_3_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_3_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_3_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_3_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_4_clock; // @[issue-unit.scala 157:73]
  wire  slots_4_reset; // @[issue-unit.scala 157:73]
  wire  slots_4_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_request; // @[issue-unit.scala 157:73]
  wire  slots_4_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_4_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_4_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_4_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_4_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_4_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_5_clock; // @[issue-unit.scala 157:73]
  wire  slots_5_reset; // @[issue-unit.scala 157:73]
  wire  slots_5_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_request; // @[issue-unit.scala 157:73]
  wire  slots_5_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_5_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_5_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_5_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_5_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_5_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_6_clock; // @[issue-unit.scala 157:73]
  wire  slots_6_reset; // @[issue-unit.scala 157:73]
  wire  slots_6_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_request; // @[issue-unit.scala 157:73]
  wire  slots_6_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_6_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_6_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_6_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_6_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_6_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_7_clock; // @[issue-unit.scala 157:73]
  wire  slots_7_reset; // @[issue-unit.scala 157:73]
  wire  slots_7_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_request; // @[issue-unit.scala 157:73]
  wire  slots_7_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_7_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_7_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_7_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_7_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_7_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_8_clock; // @[issue-unit.scala 157:73]
  wire  slots_8_reset; // @[issue-unit.scala 157:73]
  wire  slots_8_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_request; // @[issue-unit.scala 157:73]
  wire  slots_8_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_8_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_8_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_8_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_8_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_8_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_9_clock; // @[issue-unit.scala 157:73]
  wire  slots_9_reset; // @[issue-unit.scala 157:73]
  wire  slots_9_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_request; // @[issue-unit.scala 157:73]
  wire  slots_9_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_9_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_9_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_9_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_9_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_9_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_10_clock; // @[issue-unit.scala 157:73]
  wire  slots_10_reset; // @[issue-unit.scala 157:73]
  wire  slots_10_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_request; // @[issue-unit.scala 157:73]
  wire  slots_10_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_10_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_10_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_10_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_10_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_10_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_11_clock; // @[issue-unit.scala 157:73]
  wire  slots_11_reset; // @[issue-unit.scala 157:73]
  wire  slots_11_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_request; // @[issue-unit.scala 157:73]
  wire  slots_11_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_11_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_11_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_11_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_11_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_11_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_12_clock; // @[issue-unit.scala 157:73]
  wire  slots_12_reset; // @[issue-unit.scala 157:73]
  wire  slots_12_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_request; // @[issue-unit.scala 157:73]
  wire  slots_12_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_12_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_12_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_12_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_12_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_12_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_13_clock; // @[issue-unit.scala 157:73]
  wire  slots_13_reset; // @[issue-unit.scala 157:73]
  wire  slots_13_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_request; // @[issue-unit.scala 157:73]
  wire  slots_13_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_13_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_13_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_13_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_13_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_13_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_14_clock; // @[issue-unit.scala 157:73]
  wire  slots_14_reset; // @[issue-unit.scala 157:73]
  wire  slots_14_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_request; // @[issue-unit.scala 157:73]
  wire  slots_14_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_14_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_14_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_14_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_14_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_14_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_15_clock; // @[issue-unit.scala 157:73]
  wire  slots_15_reset; // @[issue-unit.scala 157:73]
  wire  slots_15_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_request; // @[issue-unit.scala 157:73]
  wire  slots_15_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_15_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_15_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_15_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_15_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_15_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_16_clock; // @[issue-unit.scala 157:73]
  wire  slots_16_reset; // @[issue-unit.scala 157:73]
  wire  slots_16_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_request; // @[issue-unit.scala 157:73]
  wire  slots_16_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_16_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_16_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_16_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_16_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_16_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_16_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_16_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_16_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_16_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_16_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_16_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_16_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_16_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_16_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_16_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_16_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_16_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_16_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_16_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_16_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_16_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_16_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_16_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_16_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_16_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_16_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_16_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_16_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_16_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_16_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_16_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_16_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_16_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_16_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_16_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_16_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_17_clock; // @[issue-unit.scala 157:73]
  wire  slots_17_reset; // @[issue-unit.scala 157:73]
  wire  slots_17_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_request; // @[issue-unit.scala 157:73]
  wire  slots_17_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_17_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_17_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_17_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_17_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_17_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_17_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_17_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_17_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_17_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_17_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_17_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_17_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_17_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_17_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_17_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_17_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_17_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_17_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_17_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_17_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_17_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_17_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_17_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_17_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_17_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_17_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_17_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_17_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_17_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_17_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_17_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_17_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_17_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_17_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_17_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_17_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_18_clock; // @[issue-unit.scala 157:73]
  wire  slots_18_reset; // @[issue-unit.scala 157:73]
  wire  slots_18_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_request; // @[issue-unit.scala 157:73]
  wire  slots_18_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_18_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_18_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_18_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_18_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_18_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_18_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_18_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_18_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_18_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_18_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_18_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_18_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_18_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_18_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_18_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_18_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_18_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_18_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_18_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_18_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_18_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_18_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_18_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_18_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_18_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_18_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_18_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_18_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_18_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_18_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_18_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_18_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_18_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_18_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_18_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_18_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_19_clock; // @[issue-unit.scala 157:73]
  wire  slots_19_reset; // @[issue-unit.scala 157:73]
  wire  slots_19_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_request; // @[issue-unit.scala 157:73]
  wire  slots_19_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_19_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_19_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_19_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_19_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_19_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_19_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_19_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_19_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_19_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_19_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_2_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_3_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_4_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_19_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_19_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_19_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_19_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_19_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_19_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_19_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_19_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_19_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_19_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_19_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_19_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_19_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_19_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_19_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_19_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_19_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_19_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_19_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_19_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_19_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_19_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_19_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_19_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_19_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_19_io_debug_state; // @[issue-unit.scala 157:73]
  wire  _T = io_dis_uops_0_bits_uopc == 7'h2; // @[issue-unit.scala 131:39]
  wire  _T_3 = io_dis_uops_0_bits_uopc == 7'h43; // @[issue-unit.scala 132:39]
  wire  _T_4 = io_dis_uops_0_bits_uopc == 7'h2 & io_dis_uops_0_bits_lrs2_rtype == 2'h0 | _T_3; // @[issue-unit.scala 131:96]
  wire [1:0] _GEN_0 = _T & io_dis_uops_0_bits_lrs2_rtype != 2'h0 ? 2'h2 : io_dis_uops_0_bits_lrs2_rtype; // @[issue-unit.scala 135:102 issue-unit.scala 136:32 issue-unit.scala 124:17]
  wire  _GEN_1 = _T & io_dis_uops_0_bits_lrs2_rtype != 2'h0 ? 1'h0 : io_dis_uops_0_bits_prs2_busy; // @[issue-unit.scala 135:102 issue-unit.scala 137:32 issue-unit.scala 124:17]
  wire [1:0] uops_20_iw_state = _T_4 ? 2'h2 : 2'h1; // @[issue-unit.scala 132:54 issue-unit.scala 133:30 issue-unit.scala 127:26]
  wire [1:0] uops_20_lrs2_rtype = _T_4 ? io_dis_uops_0_bits_lrs2_rtype : _GEN_0; // @[issue-unit.scala 132:54 issue-unit.scala 124:17]
  wire  uops_20_prs2_busy = _T_4 ? io_dis_uops_0_bits_prs2_busy : _GEN_1; // @[issue-unit.scala 132:54 issue-unit.scala 124:17]
  wire  _T_8 = io_dis_uops_1_bits_uopc == 7'h2; // @[issue-unit.scala 131:39]
  wire  _T_11 = io_dis_uops_1_bits_uopc == 7'h43; // @[issue-unit.scala 132:39]
  wire  _T_12 = io_dis_uops_1_bits_uopc == 7'h2 & io_dis_uops_1_bits_lrs2_rtype == 2'h0 | _T_11; // @[issue-unit.scala 131:96]
  wire [1:0] _GEN_5 = _T_8 & io_dis_uops_1_bits_lrs2_rtype != 2'h0 ? 2'h2 : io_dis_uops_1_bits_lrs2_rtype; // @[issue-unit.scala 135:102 issue-unit.scala 136:32 issue-unit.scala 124:17]
  wire  _GEN_6 = _T_8 & io_dis_uops_1_bits_lrs2_rtype != 2'h0 ? 1'h0 : io_dis_uops_1_bits_prs2_busy; // @[issue-unit.scala 135:102 issue-unit.scala 137:32 issue-unit.scala 124:17]
  wire [1:0] uops_21_iw_state = _T_12 ? 2'h2 : 2'h1; // @[issue-unit.scala 132:54 issue-unit.scala 133:30 issue-unit.scala 127:26]
  wire [1:0] uops_21_lrs2_rtype = _T_12 ? io_dis_uops_1_bits_lrs2_rtype : _GEN_5; // @[issue-unit.scala 132:54 issue-unit.scala 124:17]
  wire  uops_21_prs2_busy = _T_12 ? io_dis_uops_1_bits_prs2_busy : _GEN_6; // @[issue-unit.scala 132:54 issue-unit.scala 124:17]
  wire  issue_slots_0_valid = slots_0_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_valid = slots_1_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_valid = slots_2_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_valid = slots_3_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_valid = slots_4_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_valid = slots_5_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_valid = slots_6_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_valid = slots_7_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_valid = slots_8_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_valid = slots_9_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_valid = slots_10_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_valid = slots_11_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_valid = slots_12_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_valid = slots_13_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_valid = slots_14_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_valid = slots_15_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_valid = slots_16_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_valid = slots_17_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_valid = slots_18_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_valid = slots_19_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_0_request = slots_0_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_0_uop_fu_code = slots_0_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_412 = issue_slots_0_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_413 = _T_412 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_423 = issue_slots_0_request & _T_413; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_429 = ~_T_423; // @[issue-unit-age-ordered.scala 122:28]
  wire [9:0] _T_427 = issue_slots_0_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_428 = _T_427 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_431 = issue_slots_0_request & ~_T_423 & _T_428; // @[issue-unit-age-ordered.scala 122:40]
  wire  issue_slots_0_grant = issue_slots_0_request & ~_T_423 & _T_428 | _T_423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_1_request = slots_1_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_1_uop_fu_code = slots_1_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_442 = issue_slots_1_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_443 = _T_442 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_453 = issue_slots_1_request & _T_443; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_455 = issue_slots_1_request & _T_443 & _T_429; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_457 = issue_slots_1_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_458 = _T_457 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_461 = issue_slots_1_request & ~_T_455 & _T_458; // @[issue-unit-age-ordered.scala 122:40]
  wire  issue_slots_1_grant = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) |
    _T_455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_73 = issue_slots_0_grant + issue_slots_1_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_3_request = slots_3_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_3_uop_fu_code = slots_3_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_502 = issue_slots_3_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_503 = _T_502 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_513 = issue_slots_3_request & _T_503; // @[issue-unit-age-ordered.scala 129:33]
  wire  issue_slots_2_request = slots_2_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_2_uop_fu_code = slots_2_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_472 = issue_slots_2_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_473 = _T_472 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_481 = issue_slots_2_request & _T_473; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_452 = _T_453 | _T_423; // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_482 = issue_slots_2_request & _T_473 | (_T_453 | _T_423); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_515 = issue_slots_3_request & _T_503 & ~_T_482; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_517 = issue_slots_3_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_518 = _T_517 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_521 = issue_slots_3_request & ~_T_515 & _T_518; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_485 = _T_481 & ~_T_452; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_487 = issue_slots_2_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_488 = _T_487 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_496 = issue_slots_2_request & ~_T_485 & _T_488; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_467 = _T_461 | _T_431; // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_497 = issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_3_grant = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 | _T_515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_4_request = slots_4_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_4_uop_fu_code = slots_4_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_532 = issue_slots_4_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_533 = _T_532 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_543 = issue_slots_4_request & _T_533; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_512 = _T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423)); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_545 = issue_slots_4_request & _T_533 & ~_T_512; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_547 = issue_slots_4_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_548 = _T_547 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_551 = issue_slots_4_request & ~_T_545 & _T_548; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_527 = _T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431)); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_4_grant = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 | _T_545; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_75 = issue_slots_3_grant + issue_slots_4_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_2_grant = _T_496 & ~_T_467 | _T_485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _GEN_7935 = {{1'd0}, issue_slots_2_grant}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_77 = _GEN_7935 + _T_75; // @[Bitwise.scala 47:55]
  wire [2:0] _T_79 = _T_73 + _T_77[1:0]; // @[Bitwise.scala 47:55]
  wire  issue_slots_5_request = slots_5_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_5_uop_fu_code = slots_5_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_562 = issue_slots_5_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_563 = _T_562 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_573 = issue_slots_5_request & _T_563; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_542 = _T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_575 = issue_slots_5_request & _T_563 & ~_T_542; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_577 = issue_slots_5_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_578 = _T_577 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_581 = issue_slots_5_request & ~_T_575 & _T_578; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_557 = _T_551 | (_T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_5_grant = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 | _T_575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_6_request = slots_6_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_6_uop_fu_code = slots_6_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_592 = issue_slots_6_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_593 = _T_592 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_603 = issue_slots_6_request & _T_593; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_572 = _T_573 | (_T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423)))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_605 = issue_slots_6_request & _T_593 & ~_T_572; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_607 = issue_slots_6_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_608 = _T_607 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_611 = issue_slots_6_request & ~_T_605 & _T_608; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_587 = _T_581 | (_T_551 | (_T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431)))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_6_grant = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 | _T_605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_81 = issue_slots_5_grant + issue_slots_6_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_8_request = slots_8_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_8_uop_fu_code = slots_8_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_652 = issue_slots_8_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_653 = _T_652 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_663 = issue_slots_8_request & _T_653; // @[issue-unit-age-ordered.scala 129:33]
  wire  issue_slots_7_request = slots_7_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_7_uop_fu_code = slots_7_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_622 = issue_slots_7_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_623 = _T_622 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_631 = issue_slots_7_request & _T_623; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_602 = _T_603 | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_632 = issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request &
    _T_473 | (_T_453 | _T_423)))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_665 = issue_slots_8_request & _T_653 & ~_T_632; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_667 = issue_slots_8_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_668 = _T_667 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_671 = issue_slots_8_request & ~_T_665 & _T_668; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_635 = _T_631 & ~_T_602; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_637 = issue_slots_7_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_638 = _T_637 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_646 = issue_slots_7_request & ~_T_635 & _T_638; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_617 = _T_611 | (_T_581 | (_T_551 | (_T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431))))
    ); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_647 = issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (
    issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431)))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_8_grant = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 | _T_665; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_9_request = slots_9_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_9_uop_fu_code = slots_9_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_682 = issue_slots_9_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_683 = _T_682 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_693 = issue_slots_9_request & _T_683; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_662 = _T_663 | (issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (
    issue_slots_2_request & _T_473 | (_T_453 | _T_423))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_695 = issue_slots_9_request & _T_683 & ~_T_662; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_697 = issue_slots_9_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_698 = _T_697 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_701 = issue_slots_9_request & ~_T_695 & _T_698; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_677 = _T_671 | (issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (
    issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_9_grant = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 | _T_695; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_83 = issue_slots_8_grant + issue_slots_9_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_7_grant = _T_646 & ~_T_617 | _T_635; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _GEN_7936 = {{1'd0}, issue_slots_7_grant}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_85 = _GEN_7936 + _T_83; // @[Bitwise.scala 47:55]
  wire [2:0] _T_87 = _T_81 + _T_85[1:0]; // @[Bitwise.scala 47:55]
  wire [3:0] _T_89 = _T_79 + _T_87; // @[Bitwise.scala 47:55]
  wire  issue_slots_10_request = slots_10_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_10_uop_fu_code = slots_10_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_712 = issue_slots_10_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_713 = _T_712 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_723 = issue_slots_10_request & _T_713; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_692 = _T_693 | (_T_663 | (issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (
    issue_slots_2_request & _T_473 | (_T_453 | _T_423)))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_725 = issue_slots_10_request & _T_713 & ~_T_692; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_727 = issue_slots_10_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_728 = _T_727 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_731 = issue_slots_10_request & ~_T_725 & _T_728; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_707 = _T_701 | (_T_671 | (issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 |
    (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431)))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_10_grant = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 | _T_725; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_11_request = slots_11_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_11_uop_fu_code = slots_11_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_742 = issue_slots_11_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_743 = _T_742 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_753 = issue_slots_11_request & _T_743; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_722 = _T_723 | (_T_693 | (_T_663 | (issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 |
    (issue_slots_2_request & _T_473 | (_T_453 | _T_423))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_755 = issue_slots_11_request & _T_743 & ~_T_722; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_757 = issue_slots_11_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_758 = _T_757 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_761 = issue_slots_11_request & ~_T_755 & _T_758; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_737 = _T_731 | (_T_701 | (_T_671 | (issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 |
    (_T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_11_grant = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 | _T_755; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_91 = issue_slots_10_grant + issue_slots_11_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_13_request = slots_13_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_13_uop_fu_code = slots_13_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_802 = issue_slots_13_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_803 = _T_802 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_813 = issue_slots_13_request & _T_803; // @[issue-unit-age-ordered.scala 129:33]
  wire  issue_slots_12_request = slots_12_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_12_uop_fu_code = slots_12_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_772 = issue_slots_12_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_773 = _T_772 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_781 = issue_slots_12_request & _T_773; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_752 = _T_753 | (_T_723 | (_T_693 | (_T_663 | (issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 |
    (_T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423)))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_782 = issue_slots_12_request & _T_773 | (_T_753 | (_T_723 | (_T_693 | (_T_663 | (issue_slots_7_request &
    _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_815 = issue_slots_13_request & _T_803 & ~_T_782; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_817 = issue_slots_13_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_818 = _T_817 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_821 = issue_slots_13_request & ~_T_815 & _T_818; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_785 = _T_781 & ~_T_752; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_787 = issue_slots_12_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_788 = _T_787 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_796 = issue_slots_12_request & ~_T_785 & _T_788; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_767 = _T_761 | (_T_731 | (_T_701 | (_T_671 | (issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 |
    (_T_551 | (_T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431)))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_797 = issue_slots_12_request & ~_T_785 & _T_788 | (_T_761 | (_T_731 | (_T_701 | (_T_671 | (
    issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (issue_slots_2_request & ~_T_485
     & _T_488 | (_T_461 | _T_431))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_13_grant = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 | _T_815; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_14_request = slots_14_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_14_uop_fu_code = slots_14_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_832 = issue_slots_14_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_833 = _T_832 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_843 = issue_slots_14_request & _T_833; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_812 = _T_813 | (issue_slots_12_request & _T_773 | (_T_753 | (_T_723 | (_T_693 | (_T_663 | (
    issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (_T_453
     | _T_423)))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_845 = issue_slots_14_request & _T_833 & ~_T_812; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_847 = issue_slots_14_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_848 = _T_847 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_851 = issue_slots_14_request & ~_T_845 & _T_848; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_827 = _T_821 | (issue_slots_12_request & ~_T_785 & _T_788 | (_T_761 | (_T_731 | (_T_701 | (_T_671 | (
    issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (issue_slots_2_request & ~_T_485
     & _T_488 | (_T_461 | _T_431)))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_14_grant = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 | _T_845; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_93 = issue_slots_13_grant + issue_slots_14_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_12_grant = _T_796 & ~_T_767 | _T_785; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _GEN_7937 = {{1'd0}, issue_slots_12_grant}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_95 = _GEN_7937 + _T_93; // @[Bitwise.scala 47:55]
  wire [2:0] _T_97 = _T_91 + _T_95[1:0]; // @[Bitwise.scala 47:55]
  wire  issue_slots_15_request = slots_15_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_15_uop_fu_code = slots_15_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_862 = issue_slots_15_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_863 = _T_862 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_873 = issue_slots_15_request & _T_863; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_842 = _T_843 | (_T_813 | (issue_slots_12_request & _T_773 | (_T_753 | (_T_723 | (_T_693 | (_T_663 | (
    issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (_T_453
     | _T_423))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_875 = issue_slots_15_request & _T_863 & ~_T_842; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_877 = issue_slots_15_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_878 = _T_877 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_881 = issue_slots_15_request & ~_T_875 & _T_878; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_857 = _T_851 | (_T_821 | (issue_slots_12_request & ~_T_785 & _T_788 | (_T_761 | (_T_731 | (_T_701 | (_T_671
     | (issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (issue_slots_2_request & ~
    _T_485 & _T_488 | (_T_461 | _T_431))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_15_grant = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 | _T_875; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_16_request = slots_16_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_16_uop_fu_code = slots_16_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_892 = issue_slots_16_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_893 = _T_892 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_903 = issue_slots_16_request & _T_893; // @[issue-unit-age-ordered.scala 129:33]
  wire  _T_872 = _T_873 | (_T_843 | (_T_813 | (issue_slots_12_request & _T_773 | (_T_753 | (_T_723 | (_T_693 | (_T_663
     | (issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (
    _T_453 | _T_423)))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_905 = issue_slots_16_request & _T_893 & ~_T_872; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_907 = issue_slots_16_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_908 = _T_907 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_911 = issue_slots_16_request & ~_T_905 & _T_908; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_887 = _T_881 | (_T_851 | (_T_821 | (issue_slots_12_request & ~_T_785 & _T_788 | (_T_761 | (_T_731 | (_T_701
     | (_T_671 | (issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (
    issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431)))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_16_grant = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 | _T_905; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_99 = issue_slots_15_grant + issue_slots_16_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_18_request = slots_18_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_18_uop_fu_code = slots_18_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_952 = issue_slots_18_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_953 = _T_952 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_963 = issue_slots_18_request & _T_953; // @[issue-unit-age-ordered.scala 129:33]
  wire  issue_slots_17_request = slots_17_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_17_uop_fu_code = slots_17_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_922 = issue_slots_17_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_923 = _T_922 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_931 = issue_slots_17_request & _T_923; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_902 = _T_903 | (_T_873 | (_T_843 | (_T_813 | (issue_slots_12_request & _T_773 | (_T_753 | (_T_723 | (_T_693
     | (_T_663 | (issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request &
    _T_473 | (_T_453 | _T_423))))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_932 = issue_slots_17_request & _T_923 | (_T_903 | (_T_873 | (_T_843 | (_T_813 | (issue_slots_12_request &
    _T_773 | (_T_753 | (_T_723 | (_T_693 | (_T_663 | (issue_slots_7_request & _T_623 | (_T_603 | (_T_573 | (_T_543 | (
    _T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423)))))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_965 = issue_slots_18_request & _T_953 & ~_T_932; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_967 = issue_slots_18_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_968 = _T_967 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_971 = issue_slots_18_request & ~_T_965 & _T_968; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_935 = _T_931 & ~_T_902; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_937 = issue_slots_17_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_938 = _T_937 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_946 = issue_slots_17_request & ~_T_935 & _T_938; // @[issue-unit-age-ordered.scala 128:52]
  wire  _T_917 = _T_911 | (_T_881 | (_T_851 | (_T_821 | (issue_slots_12_request & ~_T_785 & _T_788 | (_T_761 | (_T_731
     | (_T_701 | (_T_671 | (issue_slots_7_request & ~_T_635 & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (
    issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431))))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_947 = issue_slots_17_request & ~_T_935 & _T_938 | (_T_911 | (_T_881 | (_T_851 | (_T_821 | (
    issue_slots_12_request & ~_T_785 & _T_788 | (_T_761 | (_T_731 | (_T_701 | (_T_671 | (issue_slots_7_request & ~_T_635
     & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431))))
    )))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_18_grant = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 | _T_965; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire  issue_slots_19_request = slots_19_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_19_uop_fu_code = slots_19_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_982 = issue_slots_19_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_983 = _T_982 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_962 = _T_963 | (issue_slots_17_request & _T_923 | (_T_903 | (_T_873 | (_T_843 | (_T_813 | (
    issue_slots_12_request & _T_773 | (_T_753 | (_T_723 | (_T_693 | (_T_663 | (issue_slots_7_request & _T_623 | (_T_603
     | (_T_573 | (_T_543 | (_T_513 | (issue_slots_2_request & _T_473 | (_T_453 | _T_423))))))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  _T_995 = issue_slots_19_request & _T_983 & ~_T_962; // @[issue-unit-age-ordered.scala 129:49]
  wire [9:0] _T_997 = issue_slots_19_uop_fu_code & io_fu_types_1; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_998 = _T_997 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_977 = _T_971 | (issue_slots_17_request & ~_T_935 & _T_938 | (_T_911 | (_T_881 | (_T_851 | (_T_821 | (
    issue_slots_12_request & ~_T_785 & _T_788 | (_T_761 | (_T_731 | (_T_701 | (_T_671 | (issue_slots_7_request & ~_T_635
     & _T_638 | (_T_611 | (_T_581 | (_T_551 | (_T_521 | (issue_slots_2_request & ~_T_485 & _T_488 | (_T_461 | _T_431))))
    ))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_19_grant = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 | _T_995; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _T_101 = issue_slots_18_grant + issue_slots_19_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_17_grant = _T_946 & ~_T_917 | _T_935; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  wire [1:0] _GEN_7938 = {{1'd0}, issue_slots_17_grant}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_103 = _GEN_7938 + _T_101; // @[Bitwise.scala 47:55]
  wire [2:0] _T_105 = _T_99 + _T_103[1:0]; // @[Bitwise.scala 47:55]
  wire [3:0] _T_107 = _T_97 + _T_105; // @[Bitwise.scala 47:55]
  wire [4:0] _T_109 = _T_89 + _T_107; // @[Bitwise.scala 47:55]
  wire  vacants_0 = ~issue_slots_0_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_1 = ~issue_slots_1_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_2 = ~issue_slots_2_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_3 = ~issue_slots_3_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_4 = ~issue_slots_4_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_5 = ~issue_slots_5_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_6 = ~issue_slots_6_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_7 = ~issue_slots_7_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_8 = ~issue_slots_8_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_9 = ~issue_slots_9_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_10 = ~issue_slots_10_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_11 = ~issue_slots_11_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_12 = ~issue_slots_12_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_13 = ~issue_slots_13_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_14 = ~issue_slots_14_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_15 = ~issue_slots_15_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_16 = ~issue_slots_16_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_17 = ~issue_slots_17_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_18 = ~issue_slots_18_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_19 = ~issue_slots_19_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_20 = ~io_dis_uops_0_valid; // @[issue-unit-age-ordered.scala 39:82]
  wire [2:0] _GEN_11 = vacants_0 ? 3'h1 : 3'h0; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_128 = {_GEN_11[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_12 = ~_GEN_11[1] & vacants_1 ? _T_128 : {{1'd0}, _GEN_11[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_13 = _GEN_11[1:0] == 2'h0 & vacants_1 ? 3'h1 : _GEN_12; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_134 = {_GEN_13[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_14 = ~_GEN_13[1] & vacants_2 ? _T_134 : {{1'd0}, _GEN_13[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_15 = _GEN_13[1:0] == 2'h0 & vacants_2 ? 3'h1 : _GEN_14; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_140 = {_GEN_15[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_16 = ~_GEN_15[1] & vacants_3 ? _T_140 : {{1'd0}, _GEN_15[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_17 = _GEN_15[1:0] == 2'h0 & vacants_3 ? 3'h1 : _GEN_16; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_146 = {_GEN_17[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_18 = ~_GEN_17[1] & vacants_4 ? _T_146 : {{1'd0}, _GEN_17[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_19 = _GEN_17[1:0] == 2'h0 & vacants_4 ? 3'h1 : _GEN_18; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_152 = {_GEN_19[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_20 = ~_GEN_19[1] & vacants_5 ? _T_152 : {{1'd0}, _GEN_19[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_21 = _GEN_19[1:0] == 2'h0 & vacants_5 ? 3'h1 : _GEN_20; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_158 = {_GEN_21[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_22 = ~_GEN_21[1] & vacants_6 ? _T_158 : {{1'd0}, _GEN_21[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_23 = _GEN_21[1:0] == 2'h0 & vacants_6 ? 3'h1 : _GEN_22; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_164 = {_GEN_23[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_24 = ~_GEN_23[1] & vacants_7 ? _T_164 : {{1'd0}, _GEN_23[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_25 = _GEN_23[1:0] == 2'h0 & vacants_7 ? 3'h1 : _GEN_24; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_170 = {_GEN_25[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_26 = ~_GEN_25[1] & vacants_8 ? _T_170 : {{1'd0}, _GEN_25[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_27 = _GEN_25[1:0] == 2'h0 & vacants_8 ? 3'h1 : _GEN_26; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_176 = {_GEN_27[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_28 = ~_GEN_27[1] & vacants_9 ? _T_176 : {{1'd0}, _GEN_27[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_29 = _GEN_27[1:0] == 2'h0 & vacants_9 ? 3'h1 : _GEN_28; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_182 = {_GEN_29[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_30 = ~_GEN_29[1] & vacants_10 ? _T_182 : {{1'd0}, _GEN_29[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_31 = _GEN_29[1:0] == 2'h0 & vacants_10 ? 3'h1 : _GEN_30; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_188 = {_GEN_31[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_32 = ~_GEN_31[1] & vacants_11 ? _T_188 : {{1'd0}, _GEN_31[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_33 = _GEN_31[1:0] == 2'h0 & vacants_11 ? 3'h1 : _GEN_32; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_194 = {_GEN_33[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_34 = ~_GEN_33[1] & vacants_12 ? _T_194 : {{1'd0}, _GEN_33[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_35 = _GEN_33[1:0] == 2'h0 & vacants_12 ? 3'h1 : _GEN_34; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_200 = {_GEN_35[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_36 = ~_GEN_35[1] & vacants_13 ? _T_200 : {{1'd0}, _GEN_35[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_37 = _GEN_35[1:0] == 2'h0 & vacants_13 ? 3'h1 : _GEN_36; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_206 = {_GEN_37[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_38 = ~_GEN_37[1] & vacants_14 ? _T_206 : {{1'd0}, _GEN_37[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_39 = _GEN_37[1:0] == 2'h0 & vacants_14 ? 3'h1 : _GEN_38; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_212 = {_GEN_39[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_40 = ~_GEN_39[1] & vacants_15 ? _T_212 : {{1'd0}, _GEN_39[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_41 = _GEN_39[1:0] == 2'h0 & vacants_15 ? 3'h1 : _GEN_40; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_218 = {_GEN_41[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_42 = ~_GEN_41[1] & vacants_16 ? _T_218 : {{1'd0}, _GEN_41[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_43 = _GEN_41[1:0] == 2'h0 & vacants_16 ? 3'h1 : _GEN_42; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_224 = {_GEN_43[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_44 = ~_GEN_43[1] & vacants_17 ? _T_224 : {{1'd0}, _GEN_43[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_45 = _GEN_43[1:0] == 2'h0 & vacants_17 ? 3'h1 : _GEN_44; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_230 = {_GEN_45[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_46 = ~_GEN_45[1] & vacants_18 ? _T_230 : {{1'd0}, _GEN_45[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_47 = _GEN_45[1:0] == 2'h0 & vacants_18 ? 3'h1 : _GEN_46; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_236 = {_GEN_47[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_48 = ~_GEN_47[1] & vacants_19 ? _T_236 : {{1'd0}, _GEN_47[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_49 = _GEN_47[1:0] == 2'h0 & vacants_19 ? 3'h1 : _GEN_48; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_242 = {_GEN_49[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_50 = ~_GEN_49[1] & vacants_20 ? _T_242 : {{1'd0}, _GEN_49[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_51 = _GEN_49[1:0] == 2'h0 & vacants_20 ? 3'h1 : _GEN_50; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire  _T_243 = ~io_dis_uops_0_bits_exception; // @[issue-unit-age-ordered.scala 62:57]
  wire  _T_244 = io_dis_uops_0_valid & _T_243; // @[issue-unit-age-ordered.scala 61:77]
  wire  _T_245 = ~io_dis_uops_0_bits_is_fence; // @[issue-unit-age-ordered.scala 63:57]
  wire  _T_246 = _T_244 & _T_245; // @[issue-unit-age-ordered.scala 62:80]
  wire  _T_247 = ~io_dis_uops_0_bits_is_fencei; // @[issue-unit-age-ordered.scala 64:57]
  wire  will_be_valid_20 = _T_246 & _T_247; // @[issue-unit-age-ordered.scala 63:79]
  wire  _T_248 = ~io_dis_uops_1_bits_exception; // @[issue-unit-age-ordered.scala 62:57]
  wire  _T_249 = io_dis_uops_1_valid & _T_248; // @[issue-unit-age-ordered.scala 61:77]
  wire  _T_250 = ~io_dis_uops_1_bits_is_fence; // @[issue-unit-age-ordered.scala 63:57]
  wire  _T_251 = _T_249 & _T_250; // @[issue-unit-age-ordered.scala 62:80]
  wire  _T_252 = ~io_dis_uops_1_bits_is_fencei; // @[issue-unit-age-ordered.scala 64:57]
  wire  will_be_valid_21 = _T_251 & _T_252; // @[issue-unit-age-ordered.scala 63:79]
  wire  issue_slots_1_will_be_valid = slots_1_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_52 = _GEN_11[1:0] == 2'h1 & issue_slots_1_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire [1:0] issue_slots_1_out_uop_debug_tsrc = slots_1_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_debug_fsrc = slots_1_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_bp_xcpt_if = slots_1_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_bp_debug_if = slots_1_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_xcpt_ma_if = slots_1_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_xcpt_ae_if = slots_1_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_xcpt_pf_if = slots_1_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_fp_single = slots_1_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_fp_val = slots_1_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_frs3_en = slots_1_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_lrs2_rtype = slots_1_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_lrs1_rtype = slots_1_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_dst_rtype = slots_1_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ldst_val = slots_1_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_lrs3 = slots_1_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_lrs2 = slots_1_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_lrs1 = slots_1_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_ldst = slots_1_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ldst_is_rs1 = slots_1_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_flush_on_commit = slots_1_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_unique = slots_1_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_sys_pc2epc = slots_1_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_uses_stq = slots_1_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_uses_ldq = slots_1_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_amo = slots_1_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_fencei = slots_1_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_fence = slots_1_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_mem_signed = slots_1_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_mem_size = slots_1_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_mem_cmd = slots_1_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_bypassable = slots_1_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_1_out_uop_exc_cause = slots_1_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_exception = slots_1_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_stale_pdst = slots_1_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ppred_busy = slots_1_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_prs3_busy = slots_1_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_prs2_busy = slots_1_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_prs1_busy = slots_1_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_ppred = slots_1_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_prs3 = slots_1_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_prs2 = slots_1_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_prs1 = slots_1_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_pdst = slots_1_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_rxq_idx = slots_1_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_stq_idx = slots_1_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_ldq_idx = slots_1_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_rob_idx = slots_1_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_1_out_uop_csr_addr = slots_1_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_1_out_uop_imm_packed = slots_1_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_taken = slots_1_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_pc_lob = slots_1_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_edge_inst = slots_1_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_ftq_idx = slots_1_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_br_tag = slots_1_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_1_out_uop_br_mask = slots_1_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_sfb = slots_1_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_jal = slots_1_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_jalr = slots_1_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_br = slots_1_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_iw_p2_poisoned = slots_1_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_iw_p1_poisoned = slots_1_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_iw_state = slots_1_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_ctrl_op3_sel = slots_1_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_is_std = slots_1_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_is_sta = slots_1_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_is_load = slots_1_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_csr_cmd = slots_1_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_fcn_dw = slots_1_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_ctrl_op_fcn = slots_1_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_imm_sel = slots_1_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_op2_sel = slots_1_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_ctrl_op1_sel = slots_1_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_ctrl_br_type = slots_1_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_1_out_uop_fu_code = slots_1_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_iq_type = slots_1_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_1_out_uop_debug_pc = slots_1_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_rvc = slots_1_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_1_out_uop_debug_inst = slots_1_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_1_out_uop_inst = slots_1_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_uopc = slots_1_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_address_num = slots_1_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_rob_inst_idx = slots_1_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_self_index = slots_1_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_split_num = slots_1_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_op2_sel = slots_1_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_op1_sel = slots_1_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_stale_pflag = slots_1_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_pflag_busy = slots_1_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_pwflag = slots_1_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_prflag = slots_1_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_wflag = slots_1_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_rflag = slots_1_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_lrs3_rtype = slots_1_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_shift = slots_1_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_unicore = slots_1_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_switch_off = slots_1_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_switch = slots_1_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_will_be_valid = slots_2_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_0_in_uop_valid = _GEN_13[1:0] == 2'h2 ? issue_slots_2_will_be_valid : _GEN_52; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_2_out_uop_debug_tsrc = slots_2_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_debug_fsrc = slots_2_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_bp_xcpt_if = slots_2_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_bp_debug_if = slots_2_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_xcpt_ma_if = slots_2_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_xcpt_ae_if = slots_2_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_xcpt_pf_if = slots_2_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_fp_single = slots_2_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_fp_val = slots_2_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_frs3_en = slots_2_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_lrs2_rtype = slots_2_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_lrs1_rtype = slots_2_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_dst_rtype = slots_2_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ldst_val = slots_2_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_lrs3 = slots_2_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_lrs2 = slots_2_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_lrs1 = slots_2_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_ldst = slots_2_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ldst_is_rs1 = slots_2_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_flush_on_commit = slots_2_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_unique = slots_2_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_sys_pc2epc = slots_2_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_uses_stq = slots_2_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_uses_ldq = slots_2_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_amo = slots_2_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_fencei = slots_2_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_fence = slots_2_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_mem_signed = slots_2_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_mem_size = slots_2_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_mem_cmd = slots_2_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_bypassable = slots_2_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_2_out_uop_exc_cause = slots_2_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_exception = slots_2_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_stale_pdst = slots_2_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ppred_busy = slots_2_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_prs3_busy = slots_2_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_prs2_busy = slots_2_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_prs1_busy = slots_2_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_ppred = slots_2_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_prs3 = slots_2_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_prs2 = slots_2_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_prs1 = slots_2_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_pdst = slots_2_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_rxq_idx = slots_2_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_stq_idx = slots_2_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_ldq_idx = slots_2_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_rob_idx = slots_2_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_2_out_uop_csr_addr = slots_2_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_2_out_uop_imm_packed = slots_2_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_taken = slots_2_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_pc_lob = slots_2_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_edge_inst = slots_2_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_ftq_idx = slots_2_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_br_tag = slots_2_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_2_out_uop_br_mask = slots_2_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_sfb = slots_2_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_jal = slots_2_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_jalr = slots_2_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_br = slots_2_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_iw_p2_poisoned = slots_2_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_iw_p1_poisoned = slots_2_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_iw_state = slots_2_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_ctrl_op3_sel = slots_2_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_is_std = slots_2_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_is_sta = slots_2_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_is_load = slots_2_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_csr_cmd = slots_2_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_fcn_dw = slots_2_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_ctrl_op_fcn = slots_2_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_imm_sel = slots_2_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_op2_sel = slots_2_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_ctrl_op1_sel = slots_2_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_ctrl_br_type = slots_2_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_2_out_uop_fu_code = slots_2_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_iq_type = slots_2_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_2_out_uop_debug_pc = slots_2_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_rvc = slots_2_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_2_out_uop_debug_inst = slots_2_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_2_out_uop_inst = slots_2_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_uopc = slots_2_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_address_num = slots_2_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_rob_inst_idx = slots_2_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_self_index = slots_2_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_split_num = slots_2_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_op2_sel = slots_2_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_op1_sel = slots_2_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_stale_pflag = slots_2_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_pflag_busy = slots_2_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_pwflag = slots_2_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_prflag = slots_2_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_wflag = slots_2_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_rflag = slots_2_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_lrs3_rtype = slots_2_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_shift = slots_2_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_unicore = slots_2_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_switch_off = slots_2_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_switch = slots_2_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_248 = _GEN_13[1:0] == 2'h1 & issue_slots_2_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_3_will_be_valid = slots_3_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_in_uop_valid = _GEN_15[1:0] == 2'h2 ? issue_slots_3_will_be_valid : _GEN_248; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_3_out_uop_debug_tsrc = slots_3_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_debug_fsrc = slots_3_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_bp_xcpt_if = slots_3_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_bp_debug_if = slots_3_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_xcpt_ma_if = slots_3_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_xcpt_ae_if = slots_3_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_xcpt_pf_if = slots_3_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_fp_single = slots_3_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_fp_val = slots_3_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_frs3_en = slots_3_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_lrs2_rtype = slots_3_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_lrs1_rtype = slots_3_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_dst_rtype = slots_3_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ldst_val = slots_3_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_lrs3 = slots_3_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_lrs2 = slots_3_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_lrs1 = slots_3_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_ldst = slots_3_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ldst_is_rs1 = slots_3_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_flush_on_commit = slots_3_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_unique = slots_3_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_sys_pc2epc = slots_3_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_uses_stq = slots_3_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_uses_ldq = slots_3_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_amo = slots_3_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_fencei = slots_3_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_fence = slots_3_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_mem_signed = slots_3_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_mem_size = slots_3_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_mem_cmd = slots_3_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_bypassable = slots_3_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_3_out_uop_exc_cause = slots_3_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_exception = slots_3_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_stale_pdst = slots_3_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ppred_busy = slots_3_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_prs3_busy = slots_3_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_prs2_busy = slots_3_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_prs1_busy = slots_3_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_ppred = slots_3_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_prs3 = slots_3_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_prs2 = slots_3_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_prs1 = slots_3_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_pdst = slots_3_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_rxq_idx = slots_3_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_stq_idx = slots_3_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_ldq_idx = slots_3_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_rob_idx = slots_3_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_3_out_uop_csr_addr = slots_3_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_3_out_uop_imm_packed = slots_3_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_taken = slots_3_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_pc_lob = slots_3_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_edge_inst = slots_3_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_ftq_idx = slots_3_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_br_tag = slots_3_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_3_out_uop_br_mask = slots_3_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_sfb = slots_3_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_jal = slots_3_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_jalr = slots_3_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_br = slots_3_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_iw_p2_poisoned = slots_3_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_iw_p1_poisoned = slots_3_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_iw_state = slots_3_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_ctrl_op3_sel = slots_3_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_is_std = slots_3_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_is_sta = slots_3_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_is_load = slots_3_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_csr_cmd = slots_3_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_fcn_dw = slots_3_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_ctrl_op_fcn = slots_3_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_imm_sel = slots_3_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_op2_sel = slots_3_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_ctrl_op1_sel = slots_3_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_ctrl_br_type = slots_3_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_3_out_uop_fu_code = slots_3_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_iq_type = slots_3_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_3_out_uop_debug_pc = slots_3_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_rvc = slots_3_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_3_out_uop_debug_inst = slots_3_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_3_out_uop_inst = slots_3_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_uopc = slots_3_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_address_num = slots_3_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_rob_inst_idx = slots_3_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_self_index = slots_3_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_split_num = slots_3_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_op2_sel = slots_3_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_op1_sel = slots_3_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_stale_pflag = slots_3_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_pflag_busy = slots_3_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_pwflag = slots_3_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_prflag = slots_3_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_wflag = slots_3_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_rflag = slots_3_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_lrs3_rtype = slots_3_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_shift = slots_3_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_unicore = slots_3_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_switch_off = slots_3_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_switch = slots_3_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_clear = _GEN_11[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_444 = _GEN_15[1:0] == 2'h1 & issue_slots_3_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_4_will_be_valid = slots_4_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_in_uop_valid = _GEN_17[1:0] == 2'h2 ? issue_slots_4_will_be_valid : _GEN_444; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_4_out_uop_debug_tsrc = slots_4_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_debug_fsrc = slots_4_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_bp_xcpt_if = slots_4_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_bp_debug_if = slots_4_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_xcpt_ma_if = slots_4_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_xcpt_ae_if = slots_4_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_xcpt_pf_if = slots_4_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_fp_single = slots_4_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_fp_val = slots_4_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_frs3_en = slots_4_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_lrs2_rtype = slots_4_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_lrs1_rtype = slots_4_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_dst_rtype = slots_4_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ldst_val = slots_4_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_lrs3 = slots_4_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_lrs2 = slots_4_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_lrs1 = slots_4_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_ldst = slots_4_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ldst_is_rs1 = slots_4_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_flush_on_commit = slots_4_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_unique = slots_4_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_sys_pc2epc = slots_4_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_uses_stq = slots_4_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_uses_ldq = slots_4_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_amo = slots_4_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_fencei = slots_4_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_fence = slots_4_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_mem_signed = slots_4_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_mem_size = slots_4_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_mem_cmd = slots_4_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_bypassable = slots_4_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_4_out_uop_exc_cause = slots_4_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_exception = slots_4_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_stale_pdst = slots_4_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ppred_busy = slots_4_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_prs3_busy = slots_4_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_prs2_busy = slots_4_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_prs1_busy = slots_4_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_ppred = slots_4_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_prs3 = slots_4_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_prs2 = slots_4_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_prs1 = slots_4_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_pdst = slots_4_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_rxq_idx = slots_4_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_stq_idx = slots_4_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_ldq_idx = slots_4_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_rob_idx = slots_4_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_4_out_uop_csr_addr = slots_4_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_4_out_uop_imm_packed = slots_4_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_taken = slots_4_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_pc_lob = slots_4_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_edge_inst = slots_4_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_ftq_idx = slots_4_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_br_tag = slots_4_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_4_out_uop_br_mask = slots_4_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_sfb = slots_4_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_jal = slots_4_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_jalr = slots_4_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_br = slots_4_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_iw_p2_poisoned = slots_4_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_iw_p1_poisoned = slots_4_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_iw_state = slots_4_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_ctrl_op3_sel = slots_4_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_is_std = slots_4_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_is_sta = slots_4_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_is_load = slots_4_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_csr_cmd = slots_4_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_fcn_dw = slots_4_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_ctrl_op_fcn = slots_4_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_imm_sel = slots_4_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_op2_sel = slots_4_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_ctrl_op1_sel = slots_4_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_ctrl_br_type = slots_4_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_4_out_uop_fu_code = slots_4_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_iq_type = slots_4_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_4_out_uop_debug_pc = slots_4_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_rvc = slots_4_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_4_out_uop_debug_inst = slots_4_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_4_out_uop_inst = slots_4_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_uopc = slots_4_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_address_num = slots_4_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_rob_inst_idx = slots_4_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_self_index = slots_4_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_split_num = slots_4_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_op2_sel = slots_4_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_op1_sel = slots_4_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_stale_pflag = slots_4_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_pflag_busy = slots_4_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_pwflag = slots_4_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_prflag = slots_4_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_wflag = slots_4_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_rflag = slots_4_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_lrs3_rtype = slots_4_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_shift = slots_4_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_unicore = slots_4_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_switch_off = slots_4_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_switch = slots_4_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_clear = _GEN_13[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_640 = _GEN_17[1:0] == 2'h1 & issue_slots_4_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_5_will_be_valid = slots_5_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_in_uop_valid = _GEN_19[1:0] == 2'h2 ? issue_slots_5_will_be_valid : _GEN_640; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_5_out_uop_debug_tsrc = slots_5_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_debug_fsrc = slots_5_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_bp_xcpt_if = slots_5_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_bp_debug_if = slots_5_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_xcpt_ma_if = slots_5_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_xcpt_ae_if = slots_5_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_xcpt_pf_if = slots_5_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_fp_single = slots_5_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_fp_val = slots_5_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_frs3_en = slots_5_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_lrs2_rtype = slots_5_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_lrs1_rtype = slots_5_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_dst_rtype = slots_5_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ldst_val = slots_5_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_lrs3 = slots_5_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_lrs2 = slots_5_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_lrs1 = slots_5_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_ldst = slots_5_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ldst_is_rs1 = slots_5_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_flush_on_commit = slots_5_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_unique = slots_5_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_sys_pc2epc = slots_5_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_uses_stq = slots_5_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_uses_ldq = slots_5_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_amo = slots_5_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_fencei = slots_5_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_fence = slots_5_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_mem_signed = slots_5_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_mem_size = slots_5_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_mem_cmd = slots_5_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_bypassable = slots_5_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_5_out_uop_exc_cause = slots_5_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_exception = slots_5_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_stale_pdst = slots_5_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ppred_busy = slots_5_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_prs3_busy = slots_5_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_prs2_busy = slots_5_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_prs1_busy = slots_5_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_ppred = slots_5_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_prs3 = slots_5_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_prs2 = slots_5_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_prs1 = slots_5_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_pdst = slots_5_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_rxq_idx = slots_5_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_stq_idx = slots_5_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_ldq_idx = slots_5_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_rob_idx = slots_5_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_5_out_uop_csr_addr = slots_5_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_5_out_uop_imm_packed = slots_5_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_taken = slots_5_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_pc_lob = slots_5_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_edge_inst = slots_5_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_ftq_idx = slots_5_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_br_tag = slots_5_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_5_out_uop_br_mask = slots_5_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_sfb = slots_5_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_jal = slots_5_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_jalr = slots_5_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_br = slots_5_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_iw_p2_poisoned = slots_5_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_iw_p1_poisoned = slots_5_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_iw_state = slots_5_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_ctrl_op3_sel = slots_5_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_is_std = slots_5_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_is_sta = slots_5_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_is_load = slots_5_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_csr_cmd = slots_5_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_fcn_dw = slots_5_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_ctrl_op_fcn = slots_5_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_imm_sel = slots_5_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_op2_sel = slots_5_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_ctrl_op1_sel = slots_5_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_ctrl_br_type = slots_5_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_5_out_uop_fu_code = slots_5_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_iq_type = slots_5_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_5_out_uop_debug_pc = slots_5_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_rvc = slots_5_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_5_out_uop_debug_inst = slots_5_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_5_out_uop_inst = slots_5_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_uopc = slots_5_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_address_num = slots_5_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_rob_inst_idx = slots_5_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_self_index = slots_5_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_split_num = slots_5_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_op2_sel = slots_5_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_op1_sel = slots_5_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_stale_pflag = slots_5_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_pflag_busy = slots_5_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_pwflag = slots_5_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_prflag = slots_5_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_wflag = slots_5_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_rflag = slots_5_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_lrs3_rtype = slots_5_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_shift = slots_5_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_unicore = slots_5_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_switch_off = slots_5_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_switch = slots_5_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_clear = _GEN_15[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_836 = _GEN_19[1:0] == 2'h1 & issue_slots_5_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_6_will_be_valid = slots_6_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_in_uop_valid = _GEN_21[1:0] == 2'h2 ? issue_slots_6_will_be_valid : _GEN_836; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_6_out_uop_debug_tsrc = slots_6_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_debug_fsrc = slots_6_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_bp_xcpt_if = slots_6_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_bp_debug_if = slots_6_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_xcpt_ma_if = slots_6_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_xcpt_ae_if = slots_6_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_xcpt_pf_if = slots_6_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_fp_single = slots_6_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_fp_val = slots_6_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_frs3_en = slots_6_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_lrs2_rtype = slots_6_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_lrs1_rtype = slots_6_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_dst_rtype = slots_6_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ldst_val = slots_6_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_lrs3 = slots_6_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_lrs2 = slots_6_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_lrs1 = slots_6_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_ldst = slots_6_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ldst_is_rs1 = slots_6_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_flush_on_commit = slots_6_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_unique = slots_6_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_sys_pc2epc = slots_6_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_uses_stq = slots_6_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_uses_ldq = slots_6_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_amo = slots_6_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_fencei = slots_6_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_fence = slots_6_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_mem_signed = slots_6_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_mem_size = slots_6_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_mem_cmd = slots_6_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_bypassable = slots_6_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_6_out_uop_exc_cause = slots_6_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_exception = slots_6_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_stale_pdst = slots_6_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ppred_busy = slots_6_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_prs3_busy = slots_6_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_prs2_busy = slots_6_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_prs1_busy = slots_6_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_ppred = slots_6_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_prs3 = slots_6_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_prs2 = slots_6_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_prs1 = slots_6_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_pdst = slots_6_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_rxq_idx = slots_6_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_stq_idx = slots_6_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_ldq_idx = slots_6_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_rob_idx = slots_6_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_6_out_uop_csr_addr = slots_6_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_6_out_uop_imm_packed = slots_6_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_taken = slots_6_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_pc_lob = slots_6_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_edge_inst = slots_6_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_ftq_idx = slots_6_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_br_tag = slots_6_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_6_out_uop_br_mask = slots_6_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_sfb = slots_6_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_jal = slots_6_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_jalr = slots_6_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_br = slots_6_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_iw_p2_poisoned = slots_6_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_iw_p1_poisoned = slots_6_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_iw_state = slots_6_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_ctrl_op3_sel = slots_6_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_is_std = slots_6_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_is_sta = slots_6_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_is_load = slots_6_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_csr_cmd = slots_6_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_fcn_dw = slots_6_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_ctrl_op_fcn = slots_6_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_imm_sel = slots_6_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_op2_sel = slots_6_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_ctrl_op1_sel = slots_6_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_ctrl_br_type = slots_6_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_6_out_uop_fu_code = slots_6_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_iq_type = slots_6_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_6_out_uop_debug_pc = slots_6_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_rvc = slots_6_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_6_out_uop_debug_inst = slots_6_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_6_out_uop_inst = slots_6_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_uopc = slots_6_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_address_num = slots_6_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_rob_inst_idx = slots_6_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_self_index = slots_6_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_split_num = slots_6_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_op2_sel = slots_6_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_op1_sel = slots_6_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_stale_pflag = slots_6_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_pflag_busy = slots_6_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_pwflag = slots_6_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_prflag = slots_6_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_wflag = slots_6_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_rflag = slots_6_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_lrs3_rtype = slots_6_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_shift = slots_6_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_unicore = slots_6_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_switch_off = slots_6_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_switch = slots_6_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_clear = _GEN_17[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1032 = _GEN_21[1:0] == 2'h1 & issue_slots_6_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_7_will_be_valid = slots_7_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_in_uop_valid = _GEN_23[1:0] == 2'h2 ? issue_slots_7_will_be_valid : _GEN_1032; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_7_out_uop_debug_tsrc = slots_7_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_debug_fsrc = slots_7_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_bp_xcpt_if = slots_7_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_bp_debug_if = slots_7_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_xcpt_ma_if = slots_7_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_xcpt_ae_if = slots_7_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_xcpt_pf_if = slots_7_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_fp_single = slots_7_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_fp_val = slots_7_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_frs3_en = slots_7_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_lrs2_rtype = slots_7_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_lrs1_rtype = slots_7_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_dst_rtype = slots_7_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ldst_val = slots_7_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_lrs3 = slots_7_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_lrs2 = slots_7_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_lrs1 = slots_7_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_ldst = slots_7_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ldst_is_rs1 = slots_7_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_flush_on_commit = slots_7_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_unique = slots_7_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_sys_pc2epc = slots_7_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_uses_stq = slots_7_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_uses_ldq = slots_7_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_amo = slots_7_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_fencei = slots_7_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_fence = slots_7_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_mem_signed = slots_7_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_mem_size = slots_7_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_mem_cmd = slots_7_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_bypassable = slots_7_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_7_out_uop_exc_cause = slots_7_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_exception = slots_7_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_stale_pdst = slots_7_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ppred_busy = slots_7_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_prs3_busy = slots_7_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_prs2_busy = slots_7_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_prs1_busy = slots_7_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_ppred = slots_7_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_prs3 = slots_7_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_prs2 = slots_7_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_prs1 = slots_7_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_pdst = slots_7_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_rxq_idx = slots_7_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_stq_idx = slots_7_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_ldq_idx = slots_7_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_rob_idx = slots_7_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_7_out_uop_csr_addr = slots_7_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_7_out_uop_imm_packed = slots_7_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_taken = slots_7_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_pc_lob = slots_7_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_edge_inst = slots_7_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_ftq_idx = slots_7_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_br_tag = slots_7_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_7_out_uop_br_mask = slots_7_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_sfb = slots_7_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_jal = slots_7_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_jalr = slots_7_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_br = slots_7_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_iw_p2_poisoned = slots_7_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_iw_p1_poisoned = slots_7_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_iw_state = slots_7_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_ctrl_op3_sel = slots_7_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_is_std = slots_7_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_is_sta = slots_7_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_is_load = slots_7_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_csr_cmd = slots_7_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_fcn_dw = slots_7_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_ctrl_op_fcn = slots_7_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_imm_sel = slots_7_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_op2_sel = slots_7_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_ctrl_op1_sel = slots_7_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_ctrl_br_type = slots_7_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_7_out_uop_fu_code = slots_7_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_iq_type = slots_7_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_7_out_uop_debug_pc = slots_7_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_rvc = slots_7_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_7_out_uop_debug_inst = slots_7_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_7_out_uop_inst = slots_7_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_uopc = slots_7_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_address_num = slots_7_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_rob_inst_idx = slots_7_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_self_index = slots_7_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_split_num = slots_7_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_op2_sel = slots_7_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_op1_sel = slots_7_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_stale_pflag = slots_7_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_pflag_busy = slots_7_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_pwflag = slots_7_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_prflag = slots_7_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_wflag = slots_7_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_rflag = slots_7_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_lrs3_rtype = slots_7_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_shift = slots_7_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_unicore = slots_7_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_switch_off = slots_7_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_switch = slots_7_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_clear = _GEN_19[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1228 = _GEN_23[1:0] == 2'h1 & issue_slots_7_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_8_will_be_valid = slots_8_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_in_uop_valid = _GEN_25[1:0] == 2'h2 ? issue_slots_8_will_be_valid : _GEN_1228; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_8_out_uop_debug_tsrc = slots_8_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_debug_fsrc = slots_8_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_bp_xcpt_if = slots_8_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_bp_debug_if = slots_8_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_xcpt_ma_if = slots_8_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_xcpt_ae_if = slots_8_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_xcpt_pf_if = slots_8_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_fp_single = slots_8_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_fp_val = slots_8_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_frs3_en = slots_8_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_lrs2_rtype = slots_8_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_lrs1_rtype = slots_8_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_dst_rtype = slots_8_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ldst_val = slots_8_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_lrs3 = slots_8_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_lrs2 = slots_8_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_lrs1 = slots_8_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_ldst = slots_8_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ldst_is_rs1 = slots_8_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_flush_on_commit = slots_8_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_unique = slots_8_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_sys_pc2epc = slots_8_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_uses_stq = slots_8_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_uses_ldq = slots_8_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_amo = slots_8_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_fencei = slots_8_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_fence = slots_8_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_mem_signed = slots_8_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_mem_size = slots_8_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_mem_cmd = slots_8_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_bypassable = slots_8_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_8_out_uop_exc_cause = slots_8_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_exception = slots_8_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_stale_pdst = slots_8_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ppred_busy = slots_8_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_prs3_busy = slots_8_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_prs2_busy = slots_8_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_prs1_busy = slots_8_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_ppred = slots_8_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_prs3 = slots_8_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_prs2 = slots_8_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_prs1 = slots_8_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_pdst = slots_8_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_rxq_idx = slots_8_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_stq_idx = slots_8_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_ldq_idx = slots_8_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_rob_idx = slots_8_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_8_out_uop_csr_addr = slots_8_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_8_out_uop_imm_packed = slots_8_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_taken = slots_8_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_pc_lob = slots_8_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_edge_inst = slots_8_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_ftq_idx = slots_8_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_br_tag = slots_8_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_8_out_uop_br_mask = slots_8_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_sfb = slots_8_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_jal = slots_8_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_jalr = slots_8_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_br = slots_8_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_iw_p2_poisoned = slots_8_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_iw_p1_poisoned = slots_8_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_iw_state = slots_8_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_ctrl_op3_sel = slots_8_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_is_std = slots_8_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_is_sta = slots_8_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_is_load = slots_8_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_csr_cmd = slots_8_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_fcn_dw = slots_8_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_ctrl_op_fcn = slots_8_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_imm_sel = slots_8_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_op2_sel = slots_8_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_ctrl_op1_sel = slots_8_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_ctrl_br_type = slots_8_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_8_out_uop_fu_code = slots_8_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_iq_type = slots_8_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_8_out_uop_debug_pc = slots_8_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_rvc = slots_8_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_8_out_uop_debug_inst = slots_8_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_8_out_uop_inst = slots_8_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_uopc = slots_8_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_address_num = slots_8_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_rob_inst_idx = slots_8_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_self_index = slots_8_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_split_num = slots_8_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_op2_sel = slots_8_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_op1_sel = slots_8_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_stale_pflag = slots_8_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_pflag_busy = slots_8_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_pwflag = slots_8_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_prflag = slots_8_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_wflag = slots_8_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_rflag = slots_8_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_lrs3_rtype = slots_8_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_shift = slots_8_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_unicore = slots_8_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_switch_off = slots_8_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_switch = slots_8_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_clear = _GEN_21[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1424 = _GEN_25[1:0] == 2'h1 & issue_slots_8_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_9_will_be_valid = slots_9_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_in_uop_valid = _GEN_27[1:0] == 2'h2 ? issue_slots_9_will_be_valid : _GEN_1424; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_9_out_uop_debug_tsrc = slots_9_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_debug_fsrc = slots_9_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_bp_xcpt_if = slots_9_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_bp_debug_if = slots_9_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_xcpt_ma_if = slots_9_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_xcpt_ae_if = slots_9_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_xcpt_pf_if = slots_9_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_fp_single = slots_9_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_fp_val = slots_9_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_frs3_en = slots_9_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_lrs2_rtype = slots_9_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_lrs1_rtype = slots_9_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_dst_rtype = slots_9_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ldst_val = slots_9_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_lrs3 = slots_9_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_lrs2 = slots_9_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_lrs1 = slots_9_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_ldst = slots_9_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ldst_is_rs1 = slots_9_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_flush_on_commit = slots_9_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_unique = slots_9_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_sys_pc2epc = slots_9_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_uses_stq = slots_9_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_uses_ldq = slots_9_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_amo = slots_9_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_fencei = slots_9_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_fence = slots_9_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_mem_signed = slots_9_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_mem_size = slots_9_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_mem_cmd = slots_9_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_bypassable = slots_9_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_9_out_uop_exc_cause = slots_9_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_exception = slots_9_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_stale_pdst = slots_9_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ppred_busy = slots_9_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_prs3_busy = slots_9_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_prs2_busy = slots_9_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_prs1_busy = slots_9_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_ppred = slots_9_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_prs3 = slots_9_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_prs2 = slots_9_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_prs1 = slots_9_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_pdst = slots_9_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_rxq_idx = slots_9_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_stq_idx = slots_9_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_ldq_idx = slots_9_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_rob_idx = slots_9_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_9_out_uop_csr_addr = slots_9_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_9_out_uop_imm_packed = slots_9_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_taken = slots_9_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_pc_lob = slots_9_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_edge_inst = slots_9_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_ftq_idx = slots_9_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_br_tag = slots_9_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_9_out_uop_br_mask = slots_9_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_sfb = slots_9_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_jal = slots_9_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_jalr = slots_9_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_br = slots_9_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_iw_p2_poisoned = slots_9_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_iw_p1_poisoned = slots_9_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_iw_state = slots_9_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_ctrl_op3_sel = slots_9_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_is_std = slots_9_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_is_sta = slots_9_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_is_load = slots_9_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_csr_cmd = slots_9_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_fcn_dw = slots_9_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_ctrl_op_fcn = slots_9_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_imm_sel = slots_9_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_op2_sel = slots_9_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_ctrl_op1_sel = slots_9_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_ctrl_br_type = slots_9_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_9_out_uop_fu_code = slots_9_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_iq_type = slots_9_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_9_out_uop_debug_pc = slots_9_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_rvc = slots_9_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_9_out_uop_debug_inst = slots_9_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_9_out_uop_inst = slots_9_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_uopc = slots_9_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_address_num = slots_9_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_rob_inst_idx = slots_9_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_self_index = slots_9_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_split_num = slots_9_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_op2_sel = slots_9_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_op1_sel = slots_9_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_stale_pflag = slots_9_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_pflag_busy = slots_9_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_pwflag = slots_9_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_prflag = slots_9_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_wflag = slots_9_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_rflag = slots_9_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_lrs3_rtype = slots_9_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_shift = slots_9_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_unicore = slots_9_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_switch_off = slots_9_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_switch = slots_9_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_clear = _GEN_23[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1620 = _GEN_27[1:0] == 2'h1 & issue_slots_9_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_10_will_be_valid = slots_10_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_in_uop_valid = _GEN_29[1:0] == 2'h2 ? issue_slots_10_will_be_valid : _GEN_1620; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_10_out_uop_debug_tsrc = slots_10_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_debug_fsrc = slots_10_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_bp_xcpt_if = slots_10_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_bp_debug_if = slots_10_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_xcpt_ma_if = slots_10_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_xcpt_ae_if = slots_10_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_xcpt_pf_if = slots_10_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_fp_single = slots_10_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_fp_val = slots_10_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_frs3_en = slots_10_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_lrs2_rtype = slots_10_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_lrs1_rtype = slots_10_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_dst_rtype = slots_10_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ldst_val = slots_10_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_lrs3 = slots_10_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_lrs2 = slots_10_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_lrs1 = slots_10_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_ldst = slots_10_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ldst_is_rs1 = slots_10_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_flush_on_commit = slots_10_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_unique = slots_10_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_sys_pc2epc = slots_10_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_uses_stq = slots_10_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_uses_ldq = slots_10_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_amo = slots_10_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_fencei = slots_10_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_fence = slots_10_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_mem_signed = slots_10_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_mem_size = slots_10_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_mem_cmd = slots_10_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_bypassable = slots_10_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_10_out_uop_exc_cause = slots_10_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_exception = slots_10_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_stale_pdst = slots_10_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ppred_busy = slots_10_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_prs3_busy = slots_10_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_prs2_busy = slots_10_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_prs1_busy = slots_10_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_ppred = slots_10_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_prs3 = slots_10_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_prs2 = slots_10_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_prs1 = slots_10_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_pdst = slots_10_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_rxq_idx = slots_10_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_stq_idx = slots_10_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_ldq_idx = slots_10_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_rob_idx = slots_10_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_10_out_uop_csr_addr = slots_10_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_10_out_uop_imm_packed = slots_10_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_taken = slots_10_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_pc_lob = slots_10_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_edge_inst = slots_10_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_ftq_idx = slots_10_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_br_tag = slots_10_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_10_out_uop_br_mask = slots_10_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_sfb = slots_10_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_jal = slots_10_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_jalr = slots_10_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_br = slots_10_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_iw_p2_poisoned = slots_10_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_iw_p1_poisoned = slots_10_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_iw_state = slots_10_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_ctrl_op3_sel = slots_10_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_is_std = slots_10_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_is_sta = slots_10_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_is_load = slots_10_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_csr_cmd = slots_10_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_fcn_dw = slots_10_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_ctrl_op_fcn = slots_10_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_imm_sel = slots_10_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_op2_sel = slots_10_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_ctrl_op1_sel = slots_10_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_ctrl_br_type = slots_10_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_10_out_uop_fu_code = slots_10_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_iq_type = slots_10_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_10_out_uop_debug_pc = slots_10_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_rvc = slots_10_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_10_out_uop_debug_inst = slots_10_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_10_out_uop_inst = slots_10_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_uopc = slots_10_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_address_num = slots_10_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_rob_inst_idx = slots_10_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_self_index = slots_10_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_split_num = slots_10_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_op2_sel = slots_10_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_op1_sel = slots_10_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_stale_pflag = slots_10_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_pflag_busy = slots_10_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_pwflag = slots_10_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_prflag = slots_10_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_wflag = slots_10_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_rflag = slots_10_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_lrs3_rtype = slots_10_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_shift = slots_10_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_unicore = slots_10_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_switch_off = slots_10_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_switch = slots_10_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_clear = _GEN_25[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1816 = _GEN_29[1:0] == 2'h1 & issue_slots_10_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_11_will_be_valid = slots_11_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_in_uop_valid = _GEN_31[1:0] == 2'h2 ? issue_slots_11_will_be_valid : _GEN_1816; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_11_out_uop_debug_tsrc = slots_11_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_debug_fsrc = slots_11_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_bp_xcpt_if = slots_11_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_bp_debug_if = slots_11_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_xcpt_ma_if = slots_11_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_xcpt_ae_if = slots_11_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_xcpt_pf_if = slots_11_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_fp_single = slots_11_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_fp_val = slots_11_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_frs3_en = slots_11_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_lrs2_rtype = slots_11_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_lrs1_rtype = slots_11_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_dst_rtype = slots_11_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ldst_val = slots_11_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_lrs3 = slots_11_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_lrs2 = slots_11_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_lrs1 = slots_11_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_ldst = slots_11_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ldst_is_rs1 = slots_11_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_flush_on_commit = slots_11_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_unique = slots_11_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_sys_pc2epc = slots_11_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_uses_stq = slots_11_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_uses_ldq = slots_11_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_amo = slots_11_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_fencei = slots_11_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_fence = slots_11_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_mem_signed = slots_11_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_mem_size = slots_11_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_mem_cmd = slots_11_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_bypassable = slots_11_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_11_out_uop_exc_cause = slots_11_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_exception = slots_11_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_stale_pdst = slots_11_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ppred_busy = slots_11_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_prs3_busy = slots_11_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_prs2_busy = slots_11_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_prs1_busy = slots_11_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_ppred = slots_11_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_prs3 = slots_11_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_prs2 = slots_11_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_prs1 = slots_11_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_pdst = slots_11_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_rxq_idx = slots_11_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_stq_idx = slots_11_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_ldq_idx = slots_11_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_rob_idx = slots_11_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_11_out_uop_csr_addr = slots_11_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_11_out_uop_imm_packed = slots_11_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_taken = slots_11_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_pc_lob = slots_11_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_edge_inst = slots_11_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_ftq_idx = slots_11_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_br_tag = slots_11_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_11_out_uop_br_mask = slots_11_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_sfb = slots_11_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_jal = slots_11_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_jalr = slots_11_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_br = slots_11_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_iw_p2_poisoned = slots_11_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_iw_p1_poisoned = slots_11_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_iw_state = slots_11_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_ctrl_op3_sel = slots_11_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_is_std = slots_11_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_is_sta = slots_11_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_is_load = slots_11_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_csr_cmd = slots_11_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_fcn_dw = slots_11_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_ctrl_op_fcn = slots_11_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_imm_sel = slots_11_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_op2_sel = slots_11_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_ctrl_op1_sel = slots_11_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_ctrl_br_type = slots_11_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_11_out_uop_fu_code = slots_11_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_iq_type = slots_11_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_11_out_uop_debug_pc = slots_11_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_rvc = slots_11_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_11_out_uop_debug_inst = slots_11_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_11_out_uop_inst = slots_11_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_uopc = slots_11_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_address_num = slots_11_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_rob_inst_idx = slots_11_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_self_index = slots_11_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_split_num = slots_11_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_op2_sel = slots_11_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_op1_sel = slots_11_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_stale_pflag = slots_11_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_pflag_busy = slots_11_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_pwflag = slots_11_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_prflag = slots_11_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_wflag = slots_11_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_rflag = slots_11_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_lrs3_rtype = slots_11_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_shift = slots_11_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_unicore = slots_11_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_switch_off = slots_11_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_switch = slots_11_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_clear = _GEN_27[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2012 = _GEN_31[1:0] == 2'h1 & issue_slots_11_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_12_will_be_valid = slots_12_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_in_uop_valid = _GEN_33[1:0] == 2'h2 ? issue_slots_12_will_be_valid : _GEN_2012; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_12_out_uop_debug_tsrc = slots_12_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_debug_fsrc = slots_12_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_bp_xcpt_if = slots_12_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_bp_debug_if = slots_12_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_xcpt_ma_if = slots_12_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_xcpt_ae_if = slots_12_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_xcpt_pf_if = slots_12_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_fp_single = slots_12_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_fp_val = slots_12_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_frs3_en = slots_12_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_lrs2_rtype = slots_12_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_lrs1_rtype = slots_12_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_dst_rtype = slots_12_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ldst_val = slots_12_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_lrs3 = slots_12_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_lrs2 = slots_12_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_lrs1 = slots_12_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_ldst = slots_12_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ldst_is_rs1 = slots_12_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_flush_on_commit = slots_12_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_unique = slots_12_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_sys_pc2epc = slots_12_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_uses_stq = slots_12_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_uses_ldq = slots_12_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_amo = slots_12_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_fencei = slots_12_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_fence = slots_12_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_mem_signed = slots_12_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_mem_size = slots_12_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_mem_cmd = slots_12_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_bypassable = slots_12_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_12_out_uop_exc_cause = slots_12_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_exception = slots_12_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_stale_pdst = slots_12_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ppred_busy = slots_12_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_prs3_busy = slots_12_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_prs2_busy = slots_12_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_prs1_busy = slots_12_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_ppred = slots_12_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_prs3 = slots_12_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_prs2 = slots_12_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_prs1 = slots_12_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_pdst = slots_12_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_rxq_idx = slots_12_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_stq_idx = slots_12_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_ldq_idx = slots_12_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_rob_idx = slots_12_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_12_out_uop_csr_addr = slots_12_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_12_out_uop_imm_packed = slots_12_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_taken = slots_12_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_pc_lob = slots_12_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_edge_inst = slots_12_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_ftq_idx = slots_12_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_br_tag = slots_12_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_12_out_uop_br_mask = slots_12_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_sfb = slots_12_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_jal = slots_12_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_jalr = slots_12_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_br = slots_12_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_iw_p2_poisoned = slots_12_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_iw_p1_poisoned = slots_12_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_iw_state = slots_12_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_ctrl_op3_sel = slots_12_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_is_std = slots_12_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_is_sta = slots_12_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_is_load = slots_12_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_ctrl_csr_cmd = slots_12_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_fcn_dw = slots_12_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_ctrl_op_fcn = slots_12_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_ctrl_imm_sel = slots_12_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_ctrl_op2_sel = slots_12_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_ctrl_op1_sel = slots_12_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_ctrl_br_type = slots_12_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_12_out_uop_fu_code = slots_12_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_iq_type = slots_12_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_12_out_uop_debug_pc = slots_12_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_rvc = slots_12_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_12_out_uop_debug_inst = slots_12_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_12_out_uop_inst = slots_12_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_uopc = slots_12_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_address_num = slots_12_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_rob_inst_idx = slots_12_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_self_index = slots_12_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_split_num = slots_12_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_op2_sel = slots_12_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_op1_sel = slots_12_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_stale_pflag = slots_12_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_pflag_busy = slots_12_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_pwflag = slots_12_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_prflag = slots_12_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_wflag = slots_12_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_rflag = slots_12_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_lrs3_rtype = slots_12_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_shift = slots_12_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_unicore = slots_12_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_switch_off = slots_12_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_switch = slots_12_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_clear = _GEN_29[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2208 = _GEN_33[1:0] == 2'h1 & issue_slots_12_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_13_will_be_valid = slots_13_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_in_uop_valid = _GEN_35[1:0] == 2'h2 ? issue_slots_13_will_be_valid : _GEN_2208; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_13_out_uop_debug_tsrc = slots_13_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_debug_fsrc = slots_13_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_bp_xcpt_if = slots_13_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_bp_debug_if = slots_13_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_xcpt_ma_if = slots_13_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_xcpt_ae_if = slots_13_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_xcpt_pf_if = slots_13_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_fp_single = slots_13_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_fp_val = slots_13_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_frs3_en = slots_13_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_lrs2_rtype = slots_13_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_lrs1_rtype = slots_13_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_dst_rtype = slots_13_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ldst_val = slots_13_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_lrs3 = slots_13_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_lrs2 = slots_13_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_lrs1 = slots_13_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_ldst = slots_13_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ldst_is_rs1 = slots_13_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_flush_on_commit = slots_13_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_unique = slots_13_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_sys_pc2epc = slots_13_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_uses_stq = slots_13_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_uses_ldq = slots_13_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_amo = slots_13_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_fencei = slots_13_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_fence = slots_13_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_mem_signed = slots_13_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_mem_size = slots_13_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_mem_cmd = slots_13_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_bypassable = slots_13_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_13_out_uop_exc_cause = slots_13_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_exception = slots_13_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_stale_pdst = slots_13_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ppred_busy = slots_13_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_prs3_busy = slots_13_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_prs2_busy = slots_13_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_prs1_busy = slots_13_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_ppred = slots_13_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_prs3 = slots_13_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_prs2 = slots_13_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_prs1 = slots_13_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_pdst = slots_13_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_rxq_idx = slots_13_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_stq_idx = slots_13_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_ldq_idx = slots_13_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_rob_idx = slots_13_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_13_out_uop_csr_addr = slots_13_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_13_out_uop_imm_packed = slots_13_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_taken = slots_13_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_pc_lob = slots_13_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_edge_inst = slots_13_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_ftq_idx = slots_13_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_br_tag = slots_13_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_13_out_uop_br_mask = slots_13_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_sfb = slots_13_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_jal = slots_13_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_jalr = slots_13_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_br = slots_13_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_iw_p2_poisoned = slots_13_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_iw_p1_poisoned = slots_13_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_iw_state = slots_13_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_ctrl_op3_sel = slots_13_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_is_std = slots_13_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_is_sta = slots_13_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_is_load = slots_13_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_ctrl_csr_cmd = slots_13_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_fcn_dw = slots_13_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_ctrl_op_fcn = slots_13_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_ctrl_imm_sel = slots_13_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_ctrl_op2_sel = slots_13_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_ctrl_op1_sel = slots_13_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_ctrl_br_type = slots_13_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_13_out_uop_fu_code = slots_13_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_iq_type = slots_13_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_13_out_uop_debug_pc = slots_13_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_rvc = slots_13_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_13_out_uop_debug_inst = slots_13_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_13_out_uop_inst = slots_13_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_uopc = slots_13_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_address_num = slots_13_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_rob_inst_idx = slots_13_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_self_index = slots_13_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_split_num = slots_13_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_op2_sel = slots_13_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_op1_sel = slots_13_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_stale_pflag = slots_13_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_pflag_busy = slots_13_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_pwflag = slots_13_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_prflag = slots_13_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_wflag = slots_13_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_rflag = slots_13_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_lrs3_rtype = slots_13_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_shift = slots_13_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_unicore = slots_13_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_switch_off = slots_13_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_switch = slots_13_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_clear = _GEN_31[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2404 = _GEN_35[1:0] == 2'h1 & issue_slots_13_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_14_will_be_valid = slots_14_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_in_uop_valid = _GEN_37[1:0] == 2'h2 ? issue_slots_14_will_be_valid : _GEN_2404; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_14_out_uop_debug_tsrc = slots_14_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_debug_fsrc = slots_14_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_bp_xcpt_if = slots_14_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_bp_debug_if = slots_14_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_xcpt_ma_if = slots_14_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_xcpt_ae_if = slots_14_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_xcpt_pf_if = slots_14_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_fp_single = slots_14_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_fp_val = slots_14_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_frs3_en = slots_14_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_lrs2_rtype = slots_14_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_lrs1_rtype = slots_14_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_dst_rtype = slots_14_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ldst_val = slots_14_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_lrs3 = slots_14_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_lrs2 = slots_14_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_lrs1 = slots_14_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_ldst = slots_14_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ldst_is_rs1 = slots_14_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_flush_on_commit = slots_14_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_unique = slots_14_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_sys_pc2epc = slots_14_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_uses_stq = slots_14_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_uses_ldq = slots_14_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_amo = slots_14_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_fencei = slots_14_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_fence = slots_14_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_mem_signed = slots_14_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_mem_size = slots_14_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_mem_cmd = slots_14_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_bypassable = slots_14_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_14_out_uop_exc_cause = slots_14_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_exception = slots_14_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_stale_pdst = slots_14_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ppred_busy = slots_14_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_prs3_busy = slots_14_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_prs2_busy = slots_14_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_prs1_busy = slots_14_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_ppred = slots_14_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_prs3 = slots_14_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_prs2 = slots_14_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_prs1 = slots_14_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_pdst = slots_14_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_rxq_idx = slots_14_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_stq_idx = slots_14_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_ldq_idx = slots_14_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_rob_idx = slots_14_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_14_out_uop_csr_addr = slots_14_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_14_out_uop_imm_packed = slots_14_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_taken = slots_14_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_pc_lob = slots_14_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_edge_inst = slots_14_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_ftq_idx = slots_14_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_br_tag = slots_14_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_14_out_uop_br_mask = slots_14_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_sfb = slots_14_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_jal = slots_14_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_jalr = slots_14_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_br = slots_14_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_iw_p2_poisoned = slots_14_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_iw_p1_poisoned = slots_14_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_iw_state = slots_14_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_ctrl_op3_sel = slots_14_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_is_std = slots_14_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_is_sta = slots_14_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_is_load = slots_14_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_ctrl_csr_cmd = slots_14_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_fcn_dw = slots_14_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_ctrl_op_fcn = slots_14_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_ctrl_imm_sel = slots_14_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_ctrl_op2_sel = slots_14_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_ctrl_op1_sel = slots_14_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_ctrl_br_type = slots_14_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_14_out_uop_fu_code = slots_14_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_iq_type = slots_14_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_14_out_uop_debug_pc = slots_14_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_rvc = slots_14_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_14_out_uop_debug_inst = slots_14_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_14_out_uop_inst = slots_14_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_uopc = slots_14_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_address_num = slots_14_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_rob_inst_idx = slots_14_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_self_index = slots_14_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_split_num = slots_14_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_op2_sel = slots_14_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_op1_sel = slots_14_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_stale_pflag = slots_14_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_pflag_busy = slots_14_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_pwflag = slots_14_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_prflag = slots_14_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_wflag = slots_14_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_rflag = slots_14_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_lrs3_rtype = slots_14_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_shift = slots_14_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_unicore = slots_14_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_switch_off = slots_14_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_switch = slots_14_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_clear = _GEN_33[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2600 = _GEN_37[1:0] == 2'h1 & issue_slots_14_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_15_will_be_valid = slots_15_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_in_uop_valid = _GEN_39[1:0] == 2'h2 ? issue_slots_15_will_be_valid : _GEN_2600; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_15_out_uop_debug_tsrc = slots_15_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_debug_fsrc = slots_15_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_bp_xcpt_if = slots_15_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_bp_debug_if = slots_15_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_xcpt_ma_if = slots_15_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_xcpt_ae_if = slots_15_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_xcpt_pf_if = slots_15_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_fp_single = slots_15_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_fp_val = slots_15_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_frs3_en = slots_15_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_lrs2_rtype = slots_15_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_lrs1_rtype = slots_15_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_dst_rtype = slots_15_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ldst_val = slots_15_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_lrs3 = slots_15_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_lrs2 = slots_15_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_lrs1 = slots_15_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_ldst = slots_15_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ldst_is_rs1 = slots_15_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_flush_on_commit = slots_15_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_unique = slots_15_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_sys_pc2epc = slots_15_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_uses_stq = slots_15_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_uses_ldq = slots_15_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_amo = slots_15_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_fencei = slots_15_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_fence = slots_15_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_mem_signed = slots_15_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_mem_size = slots_15_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_mem_cmd = slots_15_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_bypassable = slots_15_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_15_out_uop_exc_cause = slots_15_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_exception = slots_15_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_stale_pdst = slots_15_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ppred_busy = slots_15_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_prs3_busy = slots_15_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_prs2_busy = slots_15_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_prs1_busy = slots_15_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_ppred = slots_15_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_prs3 = slots_15_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_prs2 = slots_15_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_prs1 = slots_15_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_pdst = slots_15_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_rxq_idx = slots_15_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_stq_idx = slots_15_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_ldq_idx = slots_15_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_rob_idx = slots_15_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_15_out_uop_csr_addr = slots_15_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_15_out_uop_imm_packed = slots_15_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_taken = slots_15_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_pc_lob = slots_15_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_edge_inst = slots_15_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_ftq_idx = slots_15_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_br_tag = slots_15_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_15_out_uop_br_mask = slots_15_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_sfb = slots_15_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_jal = slots_15_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_jalr = slots_15_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_br = slots_15_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_iw_p2_poisoned = slots_15_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_iw_p1_poisoned = slots_15_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_iw_state = slots_15_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_ctrl_op3_sel = slots_15_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_is_std = slots_15_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_is_sta = slots_15_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_is_load = slots_15_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_ctrl_csr_cmd = slots_15_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_fcn_dw = slots_15_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_ctrl_op_fcn = slots_15_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_ctrl_imm_sel = slots_15_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_ctrl_op2_sel = slots_15_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_ctrl_op1_sel = slots_15_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_ctrl_br_type = slots_15_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_15_out_uop_fu_code = slots_15_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_iq_type = slots_15_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_15_out_uop_debug_pc = slots_15_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_rvc = slots_15_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_15_out_uop_debug_inst = slots_15_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_15_out_uop_inst = slots_15_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_uopc = slots_15_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_address_num = slots_15_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_rob_inst_idx = slots_15_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_self_index = slots_15_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_split_num = slots_15_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_op2_sel = slots_15_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_op1_sel = slots_15_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_stale_pflag = slots_15_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_pflag_busy = slots_15_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_pwflag = slots_15_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_prflag = slots_15_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_wflag = slots_15_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_rflag = slots_15_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_lrs3_rtype = slots_15_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_shift = slots_15_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_unicore = slots_15_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_switch_off = slots_15_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_switch = slots_15_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_clear = _GEN_35[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2796 = _GEN_39[1:0] == 2'h1 & issue_slots_15_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_16_will_be_valid = slots_16_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_in_uop_valid = _GEN_41[1:0] == 2'h2 ? issue_slots_16_will_be_valid : _GEN_2796; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_16_out_uop_debug_tsrc = slots_16_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_debug_fsrc = slots_16_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_bp_xcpt_if = slots_16_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_bp_debug_if = slots_16_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_xcpt_ma_if = slots_16_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_xcpt_ae_if = slots_16_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_xcpt_pf_if = slots_16_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_fp_single = slots_16_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_fp_val = slots_16_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_frs3_en = slots_16_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_lrs2_rtype = slots_16_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_lrs1_rtype = slots_16_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_dst_rtype = slots_16_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_ldst_val = slots_16_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_lrs3 = slots_16_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_lrs2 = slots_16_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_lrs1 = slots_16_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_ldst = slots_16_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_ldst_is_rs1 = slots_16_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_flush_on_commit = slots_16_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_unique = slots_16_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_sys_pc2epc = slots_16_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_uses_stq = slots_16_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_uses_ldq = slots_16_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_amo = slots_16_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_fencei = slots_16_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_fence = slots_16_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_mem_signed = slots_16_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_mem_size = slots_16_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_16_out_uop_mem_cmd = slots_16_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_bypassable = slots_16_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_16_out_uop_exc_cause = slots_16_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_exception = slots_16_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_16_out_uop_stale_pdst = slots_16_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_ppred_busy = slots_16_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_prs3_busy = slots_16_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_prs2_busy = slots_16_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_prs1_busy = slots_16_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_16_out_uop_ppred = slots_16_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_16_out_uop_prs3 = slots_16_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_16_out_uop_prs2 = slots_16_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_16_out_uop_prs1 = slots_16_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_16_out_uop_pdst = slots_16_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_rxq_idx = slots_16_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_16_out_uop_stq_idx = slots_16_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_16_out_uop_ldq_idx = slots_16_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_rob_idx = slots_16_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_16_out_uop_csr_addr = slots_16_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_16_out_uop_imm_packed = slots_16_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_taken = slots_16_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_pc_lob = slots_16_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_edge_inst = slots_16_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_16_out_uop_ftq_idx = slots_16_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_br_tag = slots_16_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_16_out_uop_br_mask = slots_16_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_sfb = slots_16_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_jal = slots_16_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_jalr = slots_16_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_br = slots_16_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_iw_p2_poisoned = slots_16_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_iw_p1_poisoned = slots_16_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_iw_state = slots_16_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_ctrl_op3_sel = slots_16_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_ctrl_is_std = slots_16_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_ctrl_is_sta = slots_16_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_ctrl_is_load = slots_16_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_16_out_uop_ctrl_csr_cmd = slots_16_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_ctrl_fcn_dw = slots_16_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_ctrl_op_fcn = slots_16_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_16_out_uop_ctrl_imm_sel = slots_16_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_16_out_uop_ctrl_op2_sel = slots_16_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_ctrl_op1_sel = slots_16_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_ctrl_br_type = slots_16_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_16_out_uop_fu_code = slots_16_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_16_out_uop_iq_type = slots_16_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_16_out_uop_debug_pc = slots_16_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_rvc = slots_16_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_16_out_uop_debug_inst = slots_16_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_16_out_uop_inst = slots_16_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_16_out_uop_uopc = slots_16_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_address_num = slots_16_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_rob_inst_idx = slots_16_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_self_index = slots_16_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_16_out_uop_split_num = slots_16_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_op2_sel = slots_16_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_op1_sel = slots_16_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_stale_pflag = slots_16_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_pflag_busy = slots_16_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_pwflag = slots_16_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_16_out_uop_prflag = slots_16_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_wflag = slots_16_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_rflag = slots_16_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_16_out_uop_lrs3_rtype = slots_16_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_16_out_uop_shift = slots_16_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_is_unicore = slots_16_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_switch_off = slots_16_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_out_uop_switch = slots_16_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_clear = _GEN_37[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2992 = _GEN_41[1:0] == 2'h1 & issue_slots_16_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_17_will_be_valid = slots_17_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_in_uop_valid = _GEN_43[1:0] == 2'h2 ? issue_slots_17_will_be_valid : _GEN_2992; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_17_out_uop_debug_tsrc = slots_17_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_debug_fsrc = slots_17_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_bp_xcpt_if = slots_17_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_bp_debug_if = slots_17_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_xcpt_ma_if = slots_17_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_xcpt_ae_if = slots_17_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_xcpt_pf_if = slots_17_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_fp_single = slots_17_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_fp_val = slots_17_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_frs3_en = slots_17_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_lrs2_rtype = slots_17_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_lrs1_rtype = slots_17_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_dst_rtype = slots_17_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_ldst_val = slots_17_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_lrs3 = slots_17_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_lrs2 = slots_17_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_lrs1 = slots_17_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_ldst = slots_17_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_ldst_is_rs1 = slots_17_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_flush_on_commit = slots_17_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_unique = slots_17_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_sys_pc2epc = slots_17_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_uses_stq = slots_17_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_uses_ldq = slots_17_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_amo = slots_17_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_fencei = slots_17_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_fence = slots_17_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_mem_signed = slots_17_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_mem_size = slots_17_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_17_out_uop_mem_cmd = slots_17_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_bypassable = slots_17_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_17_out_uop_exc_cause = slots_17_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_exception = slots_17_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_17_out_uop_stale_pdst = slots_17_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_ppred_busy = slots_17_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_prs3_busy = slots_17_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_prs2_busy = slots_17_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_prs1_busy = slots_17_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_17_out_uop_ppred = slots_17_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_17_out_uop_prs3 = slots_17_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_17_out_uop_prs2 = slots_17_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_17_out_uop_prs1 = slots_17_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_17_out_uop_pdst = slots_17_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_rxq_idx = slots_17_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_17_out_uop_stq_idx = slots_17_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_17_out_uop_ldq_idx = slots_17_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_rob_idx = slots_17_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_17_out_uop_csr_addr = slots_17_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_17_out_uop_imm_packed = slots_17_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_taken = slots_17_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_pc_lob = slots_17_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_edge_inst = slots_17_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_17_out_uop_ftq_idx = slots_17_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_br_tag = slots_17_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_17_out_uop_br_mask = slots_17_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_sfb = slots_17_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_jal = slots_17_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_jalr = slots_17_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_br = slots_17_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_iw_p2_poisoned = slots_17_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_iw_p1_poisoned = slots_17_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_iw_state = slots_17_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_ctrl_op3_sel = slots_17_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_ctrl_is_std = slots_17_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_ctrl_is_sta = slots_17_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_ctrl_is_load = slots_17_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_17_out_uop_ctrl_csr_cmd = slots_17_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_ctrl_fcn_dw = slots_17_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_ctrl_op_fcn = slots_17_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_17_out_uop_ctrl_imm_sel = slots_17_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_17_out_uop_ctrl_op2_sel = slots_17_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_ctrl_op1_sel = slots_17_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_ctrl_br_type = slots_17_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_17_out_uop_fu_code = slots_17_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_17_out_uop_iq_type = slots_17_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_17_out_uop_debug_pc = slots_17_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_rvc = slots_17_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_17_out_uop_debug_inst = slots_17_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_17_out_uop_inst = slots_17_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_17_out_uop_uopc = slots_17_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_address_num = slots_17_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_rob_inst_idx = slots_17_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_self_index = slots_17_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_17_out_uop_split_num = slots_17_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_op2_sel = slots_17_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_op1_sel = slots_17_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_stale_pflag = slots_17_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_pflag_busy = slots_17_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_pwflag = slots_17_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_17_out_uop_prflag = slots_17_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_wflag = slots_17_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_rflag = slots_17_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_17_out_uop_lrs3_rtype = slots_17_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_17_out_uop_shift = slots_17_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_is_unicore = slots_17_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_switch_off = slots_17_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_out_uop_switch = slots_17_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_clear = _GEN_39[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_3188 = _GEN_43[1:0] == 2'h1 & issue_slots_17_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_18_will_be_valid = slots_18_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_in_uop_valid = _GEN_45[1:0] == 2'h2 ? issue_slots_18_will_be_valid : _GEN_3188; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_18_out_uop_debug_tsrc = slots_18_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_debug_fsrc = slots_18_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_bp_xcpt_if = slots_18_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_bp_debug_if = slots_18_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_xcpt_ma_if = slots_18_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_xcpt_ae_if = slots_18_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_xcpt_pf_if = slots_18_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_fp_single = slots_18_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_fp_val = slots_18_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_frs3_en = slots_18_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_lrs2_rtype = slots_18_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_lrs1_rtype = slots_18_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_dst_rtype = slots_18_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_ldst_val = slots_18_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_lrs3 = slots_18_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_lrs2 = slots_18_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_lrs1 = slots_18_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_ldst = slots_18_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_ldst_is_rs1 = slots_18_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_flush_on_commit = slots_18_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_unique = slots_18_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_sys_pc2epc = slots_18_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_uses_stq = slots_18_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_uses_ldq = slots_18_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_amo = slots_18_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_fencei = slots_18_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_fence = slots_18_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_mem_signed = slots_18_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_mem_size = slots_18_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_18_out_uop_mem_cmd = slots_18_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_bypassable = slots_18_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_18_out_uop_exc_cause = slots_18_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_exception = slots_18_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_18_out_uop_stale_pdst = slots_18_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_ppred_busy = slots_18_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_prs3_busy = slots_18_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_prs2_busy = slots_18_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_prs1_busy = slots_18_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_18_out_uop_ppred = slots_18_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_18_out_uop_prs3 = slots_18_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_18_out_uop_prs2 = slots_18_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_18_out_uop_prs1 = slots_18_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_18_out_uop_pdst = slots_18_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_rxq_idx = slots_18_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_18_out_uop_stq_idx = slots_18_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_18_out_uop_ldq_idx = slots_18_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_rob_idx = slots_18_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_18_out_uop_csr_addr = slots_18_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_18_out_uop_imm_packed = slots_18_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_taken = slots_18_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_pc_lob = slots_18_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_edge_inst = slots_18_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_18_out_uop_ftq_idx = slots_18_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_br_tag = slots_18_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_18_out_uop_br_mask = slots_18_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_sfb = slots_18_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_jal = slots_18_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_jalr = slots_18_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_br = slots_18_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_iw_p2_poisoned = slots_18_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_iw_p1_poisoned = slots_18_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_iw_state = slots_18_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_ctrl_op3_sel = slots_18_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_ctrl_is_std = slots_18_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_ctrl_is_sta = slots_18_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_ctrl_is_load = slots_18_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_18_out_uop_ctrl_csr_cmd = slots_18_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_ctrl_fcn_dw = slots_18_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_ctrl_op_fcn = slots_18_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_18_out_uop_ctrl_imm_sel = slots_18_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_18_out_uop_ctrl_op2_sel = slots_18_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_ctrl_op1_sel = slots_18_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_ctrl_br_type = slots_18_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_18_out_uop_fu_code = slots_18_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_18_out_uop_iq_type = slots_18_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_18_out_uop_debug_pc = slots_18_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_rvc = slots_18_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_18_out_uop_debug_inst = slots_18_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_18_out_uop_inst = slots_18_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_18_out_uop_uopc = slots_18_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_address_num = slots_18_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_rob_inst_idx = slots_18_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_self_index = slots_18_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_18_out_uop_split_num = slots_18_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_op2_sel = slots_18_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_op1_sel = slots_18_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_stale_pflag = slots_18_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_pflag_busy = slots_18_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_pwflag = slots_18_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_18_out_uop_prflag = slots_18_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_wflag = slots_18_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_rflag = slots_18_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_18_out_uop_lrs3_rtype = slots_18_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_18_out_uop_shift = slots_18_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_is_unicore = slots_18_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_switch_off = slots_18_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_18_out_uop_switch = slots_18_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_16_clear = _GEN_41[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_3384 = _GEN_45[1:0] == 2'h1 & issue_slots_18_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_19_will_be_valid = slots_19_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_in_uop_valid = _GEN_47[1:0] == 2'h2 ? issue_slots_19_will_be_valid : _GEN_3384; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_19_out_uop_debug_tsrc = slots_19_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_debug_fsrc = slots_19_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_bp_xcpt_if = slots_19_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_bp_debug_if = slots_19_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_xcpt_ma_if = slots_19_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_xcpt_ae_if = slots_19_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_xcpt_pf_if = slots_19_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_fp_single = slots_19_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_fp_val = slots_19_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_frs3_en = slots_19_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_lrs2_rtype = slots_19_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_lrs1_rtype = slots_19_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_dst_rtype = slots_19_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_ldst_val = slots_19_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_lrs3 = slots_19_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_lrs2 = slots_19_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_lrs1 = slots_19_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_ldst = slots_19_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_ldst_is_rs1 = slots_19_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_flush_on_commit = slots_19_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_unique = slots_19_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_sys_pc2epc = slots_19_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_uses_stq = slots_19_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_uses_ldq = slots_19_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_amo = slots_19_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_fencei = slots_19_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_fence = slots_19_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_mem_signed = slots_19_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_mem_size = slots_19_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_out_uop_mem_cmd = slots_19_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_bypassable = slots_19_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_19_out_uop_exc_cause = slots_19_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_exception = slots_19_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_out_uop_stale_pdst = slots_19_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_ppred_busy = slots_19_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_prs3_busy = slots_19_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_prs2_busy = slots_19_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_prs1_busy = slots_19_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_out_uop_ppred = slots_19_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_out_uop_prs3 = slots_19_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_out_uop_prs2 = slots_19_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_out_uop_prs1 = slots_19_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_out_uop_pdst = slots_19_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_rxq_idx = slots_19_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_out_uop_stq_idx = slots_19_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_out_uop_ldq_idx = slots_19_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_rob_idx = slots_19_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_19_out_uop_csr_addr = slots_19_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_19_out_uop_imm_packed = slots_19_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_taken = slots_19_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_pc_lob = slots_19_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_edge_inst = slots_19_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_out_uop_ftq_idx = slots_19_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_br_tag = slots_19_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_19_out_uop_br_mask = slots_19_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_sfb = slots_19_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_jal = slots_19_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_jalr = slots_19_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_br = slots_19_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_iw_p2_poisoned = slots_19_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_iw_p1_poisoned = slots_19_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_iw_state = slots_19_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_ctrl_op3_sel = slots_19_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_ctrl_is_std = slots_19_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_ctrl_is_sta = slots_19_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_ctrl_is_load = slots_19_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_out_uop_ctrl_csr_cmd = slots_19_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_ctrl_fcn_dw = slots_19_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_ctrl_op_fcn = slots_19_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_out_uop_ctrl_imm_sel = slots_19_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_out_uop_ctrl_op2_sel = slots_19_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_ctrl_op1_sel = slots_19_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_ctrl_br_type = slots_19_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_19_out_uop_fu_code = slots_19_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_out_uop_iq_type = slots_19_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_19_out_uop_debug_pc = slots_19_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_rvc = slots_19_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_19_out_uop_debug_inst = slots_19_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_19_out_uop_inst = slots_19_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_out_uop_uopc = slots_19_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_address_num = slots_19_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_rob_inst_idx = slots_19_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_self_index = slots_19_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_out_uop_split_num = slots_19_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_op2_sel = slots_19_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_op1_sel = slots_19_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_stale_pflag = slots_19_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_pflag_busy = slots_19_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_pwflag = slots_19_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_out_uop_prflag = slots_19_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_wflag = slots_19_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_rflag = slots_19_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_out_uop_lrs3_rtype = slots_19_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_out_uop_shift = slots_19_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_is_unicore = slots_19_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_switch_off = slots_19_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_out_uop_switch = slots_19_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_17_clear = _GEN_43[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_3580 = _GEN_47[1:0] == 2'h1 & issue_slots_19_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_18_in_uop_valid = _GEN_49[1:0] == 2'h2 ? will_be_valid_20 : _GEN_3580; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire  issue_slots_18_clear = _GEN_45[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_3776 = _GEN_49[1:0] == 2'h1 & will_be_valid_20; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_19_in_uop_valid = _GEN_51[1:0] == 2'h2 ? will_be_valid_21 : _GEN_3776; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire  issue_slots_19_clear = _GEN_47[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  issue_slots_0_will_be_valid = slots_0_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  will_be_available_0 = ~issue_slots_0_will_be_valid & ~issue_slots_0_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_1 = (~issue_slots_1_will_be_valid | issue_slots_1_clear) & ~issue_slots_1_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_2 = (~issue_slots_2_will_be_valid | issue_slots_2_clear) & ~issue_slots_2_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_3 = (~issue_slots_3_will_be_valid | issue_slots_3_clear) & ~issue_slots_3_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_4 = (~issue_slots_4_will_be_valid | issue_slots_4_clear) & ~issue_slots_4_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_5 = (~issue_slots_5_will_be_valid | issue_slots_5_clear) & ~issue_slots_5_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_6 = (~issue_slots_6_will_be_valid | issue_slots_6_clear) & ~issue_slots_6_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_7 = (~issue_slots_7_will_be_valid | issue_slots_7_clear) & ~issue_slots_7_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_8 = (~issue_slots_8_will_be_valid | issue_slots_8_clear) & ~issue_slots_8_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_9 = (~issue_slots_9_will_be_valid | issue_slots_9_clear) & ~issue_slots_9_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_10 = (~issue_slots_10_will_be_valid | issue_slots_10_clear) & ~issue_slots_10_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_11 = (~issue_slots_11_will_be_valid | issue_slots_11_clear) & ~issue_slots_11_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_12 = (~issue_slots_12_will_be_valid | issue_slots_12_clear) & ~issue_slots_12_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_13 = (~issue_slots_13_will_be_valid | issue_slots_13_clear) & ~issue_slots_13_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_14 = (~issue_slots_14_will_be_valid | issue_slots_14_clear) & ~issue_slots_14_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_15 = (~issue_slots_15_will_be_valid | issue_slots_15_clear) & ~issue_slots_15_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_16 = (~issue_slots_16_will_be_valid | issue_slots_16_clear) & ~issue_slots_16_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_17 = (~issue_slots_17_will_be_valid | issue_slots_17_clear) & ~issue_slots_17_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_18 = (~issue_slots_18_will_be_valid | issue_slots_18_clear) & ~issue_slots_18_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_19 = (~issue_slots_19_will_be_valid | issue_slots_19_clear) & ~issue_slots_19_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire [1:0] _T_373 = will_be_available_0 + will_be_available_1; // @[Bitwise.scala 47:55]
  wire [1:0] _T_375 = will_be_available_3 + will_be_available_4; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_7939 = {{1'd0}, will_be_available_2}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_377 = _GEN_7939 + _T_375; // @[Bitwise.scala 47:55]
  wire [2:0] _T_379 = _T_373 + _T_377[1:0]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_381 = will_be_available_5 + will_be_available_6; // @[Bitwise.scala 47:55]
  wire [1:0] _T_383 = will_be_available_8 + will_be_available_9; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_7940 = {{1'd0}, will_be_available_7}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_385 = _GEN_7940 + _T_383; // @[Bitwise.scala 47:55]
  wire [2:0] _T_387 = _T_381 + _T_385[1:0]; // @[Bitwise.scala 47:55]
  wire [3:0] _T_389 = _T_379 + _T_387; // @[Bitwise.scala 47:55]
  wire [1:0] _T_391 = will_be_available_10 + will_be_available_11; // @[Bitwise.scala 47:55]
  wire [1:0] _T_393 = will_be_available_13 + will_be_available_14; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_7941 = {{1'd0}, will_be_available_12}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_395 = _GEN_7941 + _T_393; // @[Bitwise.scala 47:55]
  wire [2:0] _T_397 = _T_391 + _T_395[1:0]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_399 = will_be_available_15 + will_be_available_16; // @[Bitwise.scala 47:55]
  wire [1:0] _T_401 = will_be_available_18 + will_be_available_19; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_7942 = {{1'd0}, will_be_available_17}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_403 = _GEN_7942 + _T_401; // @[Bitwise.scala 47:55]
  wire [2:0] _T_405 = _T_399 + _T_403[1:0]; // @[Bitwise.scala 47:55]
  wire [3:0] _T_407 = _T_397 + _T_405; // @[Bitwise.scala 47:55]
  wire [4:0] num_available = _T_389 + _T_407; // @[Bitwise.scala 47:55]
  reg  REG; // @[issue-unit-age-ordered.scala 87:36]
  reg  REG_1; // @[issue-unit-age-ordered.scala 87:36]
  wire [1:0] issue_slots_0_uop_debug_tsrc = slots_0_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3973 = _T_423 ? issue_slots_0_uop_debug_tsrc : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_debug_fsrc = slots_0_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3974 = _T_423 ? issue_slots_0_uop_debug_fsrc : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bp_xcpt_if = slots_0_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3975 = _T_423 & issue_slots_0_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bp_debug_if = slots_0_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3976 = _T_423 & issue_slots_0_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_ma_if = slots_0_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3977 = _T_423 & issue_slots_0_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_ae_if = slots_0_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3978 = _T_423 & issue_slots_0_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_pf_if = slots_0_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3979 = _T_423 & issue_slots_0_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_fp_single = slots_0_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3980 = _T_423 & issue_slots_0_uop_fp_single; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_fp_val = slots_0_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3981 = _T_423 & issue_slots_0_uop_fp_val; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_frs3_en = slots_0_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3982 = _T_423 & issue_slots_0_uop_frs3_en; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_lrs2_rtype = slots_0_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3983 = _T_423 ? issue_slots_0_uop_lrs2_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 102:31]
  wire [1:0] issue_slots_0_uop_lrs1_rtype = slots_0_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3984 = _T_423 ? issue_slots_0_uop_lrs1_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 101:31]
  wire [1:0] issue_slots_0_uop_dst_rtype = slots_0_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3985 = _T_423 ? issue_slots_0_uop_dst_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ldst_val = slots_0_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3986 = _T_423 & issue_slots_0_uop_ldst_val; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs3 = slots_0_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3987 = _T_423 ? issue_slots_0_uop_lrs3 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs2 = slots_0_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3988 = _T_423 ? issue_slots_0_uop_lrs2 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs1 = slots_0_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3989 = _T_423 ? issue_slots_0_uop_lrs1 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_ldst = slots_0_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3990 = _T_423 ? issue_slots_0_uop_ldst : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ldst_is_rs1 = slots_0_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3991 = _T_423 & issue_slots_0_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_flush_on_commit = slots_0_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3992 = _T_423 & issue_slots_0_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_unique = slots_0_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3993 = _T_423 & issue_slots_0_uop_is_unique; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_sys_pc2epc = slots_0_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3994 = _T_423 & issue_slots_0_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_uses_stq = slots_0_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3995 = _T_423 & issue_slots_0_uop_uses_stq; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_uses_ldq = slots_0_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3996 = _T_423 & issue_slots_0_uop_uses_ldq; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_amo = slots_0_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3997 = _T_423 & issue_slots_0_uop_is_amo; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_fencei = slots_0_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3998 = _T_423 & issue_slots_0_uop_is_fencei; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_fence = slots_0_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3999 = _T_423 & issue_slots_0_uop_is_fence; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_mem_signed = slots_0_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4000 = _T_423 & issue_slots_0_uop_mem_signed; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_mem_size = slots_0_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4001 = _T_423 ? issue_slots_0_uop_mem_size : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_mem_cmd = slots_0_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4002 = _T_423 ? issue_slots_0_uop_mem_cmd : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bypassable = slots_0_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4003 = _T_423 & issue_slots_0_uop_bypassable; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [63:0] issue_slots_0_uop_exc_cause = slots_0_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4004 = _T_423 ? issue_slots_0_uop_exc_cause : 64'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_exception = slots_0_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4005 = _T_423 & issue_slots_0_uop_exception; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] issue_slots_0_uop_stale_pdst = slots_0_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4006 = _T_423 ? issue_slots_0_uop_stale_pdst : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ppred_busy = slots_0_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4007 = _T_423 & issue_slots_0_uop_ppred_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs3_busy = slots_0_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4008 = _T_423 & issue_slots_0_uop_prs3_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs2_busy = slots_0_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4009 = _T_423 & issue_slots_0_uop_prs2_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs1_busy = slots_0_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4010 = _T_423 & issue_slots_0_uop_prs1_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ppred = slots_0_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4011 = _T_423 ? issue_slots_0_uop_ppred : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] issue_slots_0_uop_prs3 = slots_0_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4012 = _T_423 ? issue_slots_0_uop_prs3 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 100:25]
  wire [6:0] issue_slots_0_uop_prs2 = slots_0_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4013 = _T_423 ? issue_slots_0_uop_prs2 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 99:25]
  wire [6:0] issue_slots_0_uop_prs1 = slots_0_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4014 = _T_423 ? issue_slots_0_uop_prs1 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 98:25]
  wire [6:0] issue_slots_0_uop_pdst = slots_0_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4015 = _T_423 ? issue_slots_0_uop_pdst : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_rxq_idx = slots_0_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4016 = _T_423 ? issue_slots_0_uop_rxq_idx : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_stq_idx = slots_0_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4017 = _T_423 ? issue_slots_0_uop_stq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ldq_idx = slots_0_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4018 = _T_423 ? issue_slots_0_uop_ldq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_rob_idx = slots_0_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4019 = _T_423 ? issue_slots_0_uop_rob_idx : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] issue_slots_0_uop_csr_addr = slots_0_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4020 = _T_423 ? issue_slots_0_uop_csr_addr : 12'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [19:0] issue_slots_0_uop_imm_packed = slots_0_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4021 = _T_423 ? issue_slots_0_uop_imm_packed : 20'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_taken = slots_0_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4022 = _T_423 & issue_slots_0_uop_taken; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_pc_lob = slots_0_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4023 = _T_423 ? issue_slots_0_uop_pc_lob : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_edge_inst = slots_0_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4024 = _T_423 & issue_slots_0_uop_edge_inst; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ftq_idx = slots_0_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4025 = _T_423 ? issue_slots_0_uop_ftq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_br_tag = slots_0_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4026 = _T_423 ? issue_slots_0_uop_br_tag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] issue_slots_0_uop_br_mask = slots_0_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4027 = _T_423 ? issue_slots_0_uop_br_mask : 12'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_sfb = slots_0_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4028 = _T_423 & issue_slots_0_uop_is_sfb; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_jal = slots_0_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4029 = _T_423 & issue_slots_0_uop_is_jal; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_jalr = slots_0_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4030 = _T_423 & issue_slots_0_uop_is_jalr; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_br = slots_0_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4031 = _T_423 & issue_slots_0_uop_is_br; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_iw_p2_poisoned = slots_0_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4032 = _T_423 & issue_slots_0_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_iw_p1_poisoned = slots_0_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4033 = _T_423 & issue_slots_0_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_iw_state = slots_0_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4034 = _T_423 ? issue_slots_0_uop_iw_state : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_ctrl_op3_sel = slots_0_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4035 = _T_423 ? issue_slots_0_uop_ctrl_op3_sel : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_std = slots_0_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4036 = _T_423 & issue_slots_0_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_sta = slots_0_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4037 = _T_423 & issue_slots_0_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_load = slots_0_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4038 = _T_423 & issue_slots_0_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_csr_cmd = slots_0_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4039 = _T_423 ? issue_slots_0_uop_ctrl_csr_cmd : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_fcn_dw = slots_0_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4040 = _T_423 & issue_slots_0_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_ctrl_op_fcn = slots_0_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4041 = _T_423 ? issue_slots_0_uop_ctrl_op_fcn : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_imm_sel = slots_0_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4042 = _T_423 ? issue_slots_0_uop_ctrl_imm_sel : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_op2_sel = slots_0_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4043 = _T_423 ? issue_slots_0_uop_ctrl_op2_sel : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_ctrl_op1_sel = slots_0_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4044 = _T_423 ? issue_slots_0_uop_ctrl_op1_sel : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_ctrl_br_type = slots_0_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4045 = _T_423 ? issue_slots_0_uop_ctrl_br_type : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [9:0] _GEN_4046 = _T_423 ? issue_slots_0_uop_fu_code : 10'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_iq_type = slots_0_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4047 = _T_423 ? issue_slots_0_uop_iq_type : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [39:0] issue_slots_0_uop_debug_pc = slots_0_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4048 = _T_423 ? issue_slots_0_uop_debug_pc : 40'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_rvc = slots_0_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4049 = _T_423 & issue_slots_0_uop_is_rvc; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] issue_slots_0_uop_debug_inst = slots_0_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4050 = _T_423 ? issue_slots_0_uop_debug_inst : 32'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] issue_slots_0_uop_inst = slots_0_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4051 = _T_423 ? issue_slots_0_uop_inst : 32'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] issue_slots_0_uop_uopc = slots_0_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4052 = _T_423 ? issue_slots_0_uop_uopc : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_address_num = slots_0_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4053 = _T_423 ? issue_slots_0_uop_address_num : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_rob_inst_idx = slots_0_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4054 = _T_423 ? issue_slots_0_uop_rob_inst_idx : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_self_index = slots_0_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4055 = _T_423 ? issue_slots_0_uop_self_index : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_split_num = slots_0_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4056 = _T_423 ? issue_slots_0_uop_split_num : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_op2_sel = slots_0_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4057 = _T_423 ? issue_slots_0_uop_op2_sel : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_op1_sel = slots_0_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4058 = _T_423 ? issue_slots_0_uop_op1_sel : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_stale_pflag = slots_0_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4059 = _T_423 ? issue_slots_0_uop_stale_pflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_pflag_busy = slots_0_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4060 = _T_423 & issue_slots_0_uop_pflag_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_pwflag = slots_0_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4061 = _T_423 ? issue_slots_0_uop_pwflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_prflag = slots_0_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4062 = _T_423 ? issue_slots_0_uop_prflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 105:27]
  wire  issue_slots_0_uop_wflag = slots_0_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4063 = _T_423 & issue_slots_0_uop_wflag; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_rflag = slots_0_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4064 = _T_423 & issue_slots_0_uop_rflag; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 106:26]
  wire [1:0] issue_slots_0_uop_lrs3_rtype = slots_0_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4065 = _T_423 ? issue_slots_0_uop_lrs3_rtype : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_shift = slots_0_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4066 = _T_423 ? issue_slots_0_uop_shift : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_unicore = slots_0_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4067 = _T_423 & issue_slots_0_uop_is_unicore; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_switch_off = slots_0_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4068 = _T_423 & issue_slots_0_uop_switch_off; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_switch = slots_0_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4069 = _T_423 & issue_slots_0_uop_switch; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4072 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_debug_tsrc : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4073 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_debug_fsrc : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4074 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4075 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4076 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4077 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4078 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4079 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_fp_single; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4080 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_fp_val; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4081 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_frs3_en; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4082 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_lrs2_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 102:31]
  wire [1:0] _GEN_4083 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_lrs1_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 101:31]
  wire [1:0] _GEN_4084 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_dst_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4085 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_ldst_val; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4086 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_lrs3 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4087 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_lrs2 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4088 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_lrs1 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4089 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ldst : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4090 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4091 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4092 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_unique; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4093 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4094 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_uses_stq; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4095 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_uses_ldq; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4096 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_amo; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4097 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_fencei; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4098 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_fence; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4099 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_mem_signed; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4100 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_mem_size : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] _GEN_4101 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_mem_cmd : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4102 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_bypassable; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [63:0] _GEN_4103 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_exc_cause : 64'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4104 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_exception; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] _GEN_4105 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_stale_pdst : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4106 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_ppred_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4107 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_prs3_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4108 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_prs2_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4109 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_prs1_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] _GEN_4110 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ppred : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] _GEN_4111 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_prs3 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 100:25]
  wire [6:0] _GEN_4112 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_prs2 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 99:25]
  wire [6:0] _GEN_4113 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_prs1 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 98:25]
  wire [6:0] _GEN_4114 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_pdst : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4115 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_rxq_idx : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] _GEN_4116 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_stq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] _GEN_4117 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ldq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4118 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_rob_idx : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] _GEN_4119 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_csr_addr : 12'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [19:0] _GEN_4120 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_imm_packed : 20'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4121 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_taken; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4122 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_pc_lob : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4123 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_edge_inst; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] _GEN_4124 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ftq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4125 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_br_tag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] _GEN_4126 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_br_mask : 12'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4127 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_sfb; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4128 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_jal; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4129 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_jalr; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4130 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_br; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4131 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4132 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4133 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_iw_state : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4134 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ctrl_op3_sel : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4135 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4136 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4137 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] _GEN_4138 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ctrl_csr_cmd : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4139 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4140 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ctrl_op_fcn : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] _GEN_4141 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ctrl_imm_sel : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] _GEN_4142 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ctrl_op2_sel : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] _GEN_4143 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ctrl_op1_sel : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4144 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_ctrl_br_type : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [9:0] _GEN_4145 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_fu_code : 10'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] _GEN_4146 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_iq_type : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [39:0] _GEN_4147 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_debug_pc : 40'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4148 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_rvc; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] _GEN_4149 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_debug_inst : 32'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] _GEN_4150 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_inst : 32'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] _GEN_4151 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_uopc : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4152 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_address_num : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4153 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_rob_inst_idx : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4154 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_self_index : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] _GEN_4155 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_split_num : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4156 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_op2_sel : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4157 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_op1_sel : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4158 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_stale_pflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4159 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_pflag_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4160 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_pwflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] _GEN_4161 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_prflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 105:27]
  wire  _GEN_4162 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_wflag; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4163 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_rflag; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 106:26]
  wire [1:0] _GEN_4164 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_lrs3_rtype : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] _GEN_4165 = issue_slots_0_request & ~_T_423 & _T_428 ? issue_slots_0_uop_shift : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4166 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_is_unicore; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4167 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_switch_off; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  _GEN_4168 = issue_slots_0_request & ~_T_423 & _T_428 & issue_slots_0_uop_switch; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_1_uop_debug_tsrc = slots_1_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4171 = _T_455 ? issue_slots_1_uop_debug_tsrc : _GEN_3973; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_debug_fsrc = slots_1_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4172 = _T_455 ? issue_slots_1_uop_debug_fsrc : _GEN_3974; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_bp_xcpt_if = slots_1_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4173 = _T_455 ? issue_slots_1_uop_bp_xcpt_if : _GEN_3975; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_bp_debug_if = slots_1_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4174 = _T_455 ? issue_slots_1_uop_bp_debug_if : _GEN_3976; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_xcpt_ma_if = slots_1_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4175 = _T_455 ? issue_slots_1_uop_xcpt_ma_if : _GEN_3977; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_xcpt_ae_if = slots_1_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4176 = _T_455 ? issue_slots_1_uop_xcpt_ae_if : _GEN_3978; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_xcpt_pf_if = slots_1_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4177 = _T_455 ? issue_slots_1_uop_xcpt_pf_if : _GEN_3979; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_fp_single = slots_1_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4178 = _T_455 ? issue_slots_1_uop_fp_single : _GEN_3980; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_fp_val = slots_1_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4179 = _T_455 ? issue_slots_1_uop_fp_val : _GEN_3981; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_frs3_en = slots_1_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4180 = _T_455 ? issue_slots_1_uop_frs3_en : _GEN_3982; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_lrs2_rtype = slots_1_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4181 = _T_455 ? issue_slots_1_uop_lrs2_rtype : _GEN_3983; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_lrs1_rtype = slots_1_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4182 = _T_455 ? issue_slots_1_uop_lrs1_rtype : _GEN_3984; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_dst_rtype = slots_1_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4183 = _T_455 ? issue_slots_1_uop_dst_rtype : _GEN_3985; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ldst_val = slots_1_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4184 = _T_455 ? issue_slots_1_uop_ldst_val : _GEN_3986; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_lrs3 = slots_1_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4185 = _T_455 ? issue_slots_1_uop_lrs3 : _GEN_3987; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_lrs2 = slots_1_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4186 = _T_455 ? issue_slots_1_uop_lrs2 : _GEN_3988; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_lrs1 = slots_1_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4187 = _T_455 ? issue_slots_1_uop_lrs1 : _GEN_3989; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_ldst = slots_1_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4188 = _T_455 ? issue_slots_1_uop_ldst : _GEN_3990; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ldst_is_rs1 = slots_1_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4189 = _T_455 ? issue_slots_1_uop_ldst_is_rs1 : _GEN_3991; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_flush_on_commit = slots_1_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4190 = _T_455 ? issue_slots_1_uop_flush_on_commit : _GEN_3992; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_unique = slots_1_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4191 = _T_455 ? issue_slots_1_uop_is_unique : _GEN_3993; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_sys_pc2epc = slots_1_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4192 = _T_455 ? issue_slots_1_uop_is_sys_pc2epc : _GEN_3994; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_uses_stq = slots_1_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4193 = _T_455 ? issue_slots_1_uop_uses_stq : _GEN_3995; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_uses_ldq = slots_1_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4194 = _T_455 ? issue_slots_1_uop_uses_ldq : _GEN_3996; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_amo = slots_1_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4195 = _T_455 ? issue_slots_1_uop_is_amo : _GEN_3997; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_fencei = slots_1_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4196 = _T_455 ? issue_slots_1_uop_is_fencei : _GEN_3998; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_fence = slots_1_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4197 = _T_455 ? issue_slots_1_uop_is_fence : _GEN_3999; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_mem_signed = slots_1_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4198 = _T_455 ? issue_slots_1_uop_mem_signed : _GEN_4000; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_mem_size = slots_1_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4199 = _T_455 ? issue_slots_1_uop_mem_size : _GEN_4001; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_mem_cmd = slots_1_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4200 = _T_455 ? issue_slots_1_uop_mem_cmd : _GEN_4002; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_bypassable = slots_1_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4201 = _T_455 ? issue_slots_1_uop_bypassable : _GEN_4003; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_1_uop_exc_cause = slots_1_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4202 = _T_455 ? issue_slots_1_uop_exc_cause : _GEN_4004; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_exception = slots_1_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4203 = _T_455 ? issue_slots_1_uop_exception : _GEN_4005; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_stale_pdst = slots_1_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4204 = _T_455 ? issue_slots_1_uop_stale_pdst : _GEN_4006; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ppred_busy = slots_1_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4205 = _T_455 ? issue_slots_1_uop_ppred_busy : _GEN_4007; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_prs3_busy = slots_1_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4206 = _T_455 ? issue_slots_1_uop_prs3_busy : _GEN_4008; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_prs2_busy = slots_1_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4207 = _T_455 ? issue_slots_1_uop_prs2_busy : _GEN_4009; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_prs1_busy = slots_1_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4208 = _T_455 ? issue_slots_1_uop_prs1_busy : _GEN_4010; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_ppred = slots_1_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4209 = _T_455 ? issue_slots_1_uop_ppred : _GEN_4011; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_prs3 = slots_1_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4210 = _T_455 ? issue_slots_1_uop_prs3 : _GEN_4012; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_prs2 = slots_1_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4211 = _T_455 ? issue_slots_1_uop_prs2 : _GEN_4013; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_prs1 = slots_1_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4212 = _T_455 ? issue_slots_1_uop_prs1 : _GEN_4014; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_pdst = slots_1_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4213 = _T_455 ? issue_slots_1_uop_pdst : _GEN_4015; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_rxq_idx = slots_1_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4214 = _T_455 ? issue_slots_1_uop_rxq_idx : _GEN_4016; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_stq_idx = slots_1_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4215 = _T_455 ? issue_slots_1_uop_stq_idx : _GEN_4017; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_ldq_idx = slots_1_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4216 = _T_455 ? issue_slots_1_uop_ldq_idx : _GEN_4018; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_rob_idx = slots_1_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4217 = _T_455 ? issue_slots_1_uop_rob_idx : _GEN_4019; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_1_uop_csr_addr = slots_1_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4218 = _T_455 ? issue_slots_1_uop_csr_addr : _GEN_4020; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_1_uop_imm_packed = slots_1_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4219 = _T_455 ? issue_slots_1_uop_imm_packed : _GEN_4021; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_taken = slots_1_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4220 = _T_455 ? issue_slots_1_uop_taken : _GEN_4022; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_pc_lob = slots_1_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4221 = _T_455 ? issue_slots_1_uop_pc_lob : _GEN_4023; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_edge_inst = slots_1_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4222 = _T_455 ? issue_slots_1_uop_edge_inst : _GEN_4024; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_ftq_idx = slots_1_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4223 = _T_455 ? issue_slots_1_uop_ftq_idx : _GEN_4025; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_br_tag = slots_1_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4224 = _T_455 ? issue_slots_1_uop_br_tag : _GEN_4026; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_1_uop_br_mask = slots_1_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4225 = _T_455 ? issue_slots_1_uop_br_mask : _GEN_4027; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_sfb = slots_1_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4226 = _T_455 ? issue_slots_1_uop_is_sfb : _GEN_4028; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_jal = slots_1_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4227 = _T_455 ? issue_slots_1_uop_is_jal : _GEN_4029; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_jalr = slots_1_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4228 = _T_455 ? issue_slots_1_uop_is_jalr : _GEN_4030; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_br = slots_1_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4229 = _T_455 ? issue_slots_1_uop_is_br : _GEN_4031; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_iw_p2_poisoned = slots_1_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4230 = _T_455 ? issue_slots_1_uop_iw_p2_poisoned : _GEN_4032; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_iw_p1_poisoned = slots_1_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4231 = _T_455 ? issue_slots_1_uop_iw_p1_poisoned : _GEN_4033; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_iw_state = slots_1_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4232 = _T_455 ? issue_slots_1_uop_iw_state : _GEN_4034; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_ctrl_op3_sel = slots_1_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4233 = _T_455 ? issue_slots_1_uop_ctrl_op3_sel : _GEN_4035; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_is_std = slots_1_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4234 = _T_455 ? issue_slots_1_uop_ctrl_is_std : _GEN_4036; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_is_sta = slots_1_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4235 = _T_455 ? issue_slots_1_uop_ctrl_is_sta : _GEN_4037; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_is_load = slots_1_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4236 = _T_455 ? issue_slots_1_uop_ctrl_is_load : _GEN_4038; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_ctrl_csr_cmd = slots_1_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4237 = _T_455 ? issue_slots_1_uop_ctrl_csr_cmd : _GEN_4039; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_fcn_dw = slots_1_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4238 = _T_455 ? issue_slots_1_uop_ctrl_fcn_dw : _GEN_4040; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_ctrl_op_fcn = slots_1_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4239 = _T_455 ? issue_slots_1_uop_ctrl_op_fcn : _GEN_4041; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_ctrl_imm_sel = slots_1_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4240 = _T_455 ? issue_slots_1_uop_ctrl_imm_sel : _GEN_4042; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_ctrl_op2_sel = slots_1_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4241 = _T_455 ? issue_slots_1_uop_ctrl_op2_sel : _GEN_4043; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_ctrl_op1_sel = slots_1_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4242 = _T_455 ? issue_slots_1_uop_ctrl_op1_sel : _GEN_4044; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_ctrl_br_type = slots_1_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4243 = _T_455 ? issue_slots_1_uop_ctrl_br_type : _GEN_4045; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4244 = _T_455 ? issue_slots_1_uop_fu_code : _GEN_4046; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_iq_type = slots_1_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4245 = _T_455 ? issue_slots_1_uop_iq_type : _GEN_4047; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_1_uop_debug_pc = slots_1_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4246 = _T_455 ? issue_slots_1_uop_debug_pc : _GEN_4048; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_rvc = slots_1_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4247 = _T_455 ? issue_slots_1_uop_is_rvc : _GEN_4049; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_1_uop_debug_inst = slots_1_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4248 = _T_455 ? issue_slots_1_uop_debug_inst : _GEN_4050; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_1_uop_inst = slots_1_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4249 = _T_455 ? issue_slots_1_uop_inst : _GEN_4051; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_uopc = slots_1_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4250 = _T_455 ? issue_slots_1_uop_uopc : _GEN_4052; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_address_num = slots_1_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4251 = _T_455 ? issue_slots_1_uop_address_num : _GEN_4053; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_rob_inst_idx = slots_1_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4252 = _T_455 ? issue_slots_1_uop_rob_inst_idx : _GEN_4054; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_self_index = slots_1_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4253 = _T_455 ? issue_slots_1_uop_self_index : _GEN_4055; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_split_num = slots_1_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4254 = _T_455 ? issue_slots_1_uop_split_num : _GEN_4056; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_op2_sel = slots_1_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4255 = _T_455 ? issue_slots_1_uop_op2_sel : _GEN_4057; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_op1_sel = slots_1_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4256 = _T_455 ? issue_slots_1_uop_op1_sel : _GEN_4058; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_stale_pflag = slots_1_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4257 = _T_455 ? issue_slots_1_uop_stale_pflag : _GEN_4059; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_pflag_busy = slots_1_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4258 = _T_455 ? issue_slots_1_uop_pflag_busy : _GEN_4060; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_pwflag = slots_1_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4259 = _T_455 ? issue_slots_1_uop_pwflag : _GEN_4061; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_prflag = slots_1_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4260 = _T_455 ? issue_slots_1_uop_prflag : _GEN_4062; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_wflag = slots_1_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4261 = _T_455 ? issue_slots_1_uop_wflag : _GEN_4063; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_rflag = slots_1_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4262 = _T_455 ? issue_slots_1_uop_rflag : _GEN_4064; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_lrs3_rtype = slots_1_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4263 = _T_455 ? issue_slots_1_uop_lrs3_rtype : _GEN_4065; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_shift = slots_1_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4264 = _T_455 ? issue_slots_1_uop_shift : _GEN_4066; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_unicore = slots_1_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4265 = _T_455 ? issue_slots_1_uop_is_unicore : _GEN_4067; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_switch_off = slots_1_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4266 = _T_455 ? issue_slots_1_uop_switch_off : _GEN_4068; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_switch = slots_1_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4267 = _T_455 ? issue_slots_1_uop_switch : _GEN_4069; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4270 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_debug_tsrc : _GEN_4072; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4271 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_debug_fsrc : _GEN_4073; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4272 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_bp_xcpt_if : _GEN_4074; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4273 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_bp_debug_if : _GEN_4075; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4274 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_xcpt_ma_if : _GEN_4076; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4275 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_xcpt_ae_if : _GEN_4077; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4276 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_xcpt_pf_if : _GEN_4078; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4277 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_fp_single : _GEN_4079; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4278 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_fp_val : _GEN_4080; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4279 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_frs3_en : _GEN_4081; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4280 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_lrs2_rtype : _GEN_4082; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4281 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_lrs1_rtype : _GEN_4083; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4282 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_dst_rtype : _GEN_4084; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4283 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ldst_val : _GEN_4085; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4284 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_lrs3 : _GEN_4086; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4285 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_lrs2 : _GEN_4087; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4286 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_lrs1 : _GEN_4088; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4287 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ldst : _GEN_4089; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4288 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ldst_is_rs1 : _GEN_4090; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4289 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_flush_on_commit : _GEN_4091; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4290 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_unique : _GEN_4092; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4291 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_sys_pc2epc : _GEN_4093; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4292 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_uses_stq : _GEN_4094; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4293 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_uses_ldq : _GEN_4095; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4294 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_amo : _GEN_4096; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4295 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_fencei : _GEN_4097; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4296 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_fence : _GEN_4098; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4297 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_mem_signed : _GEN_4099; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4298 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_mem_size : _GEN_4100; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4299 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_mem_cmd : _GEN_4101; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4300 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_bypassable : _GEN_4102; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_4301 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_exc_cause : _GEN_4103; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4302 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_exception : _GEN_4104; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4303 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_stale_pdst : _GEN_4105; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4304 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ppred_busy : _GEN_4106; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4305 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_prs3_busy : _GEN_4107; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4306 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_prs2_busy : _GEN_4108; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4307 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_prs1_busy : _GEN_4109; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4308 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ppred : _GEN_4110; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4309 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_prs3 : _GEN_4111; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4310 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_prs2 : _GEN_4112; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4311 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_prs1 : _GEN_4113; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4312 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_pdst : _GEN_4114; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4313 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_rxq_idx : _GEN_4115; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4314 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_stq_idx : _GEN_4116; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4315 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ldq_idx : _GEN_4117; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4316 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_rob_idx : _GEN_4118; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4317 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_csr_addr : _GEN_4119; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_4318 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_imm_packed : _GEN_4120; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4319 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_taken : _GEN_4121; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4320 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_pc_lob : _GEN_4122; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4321 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_edge_inst : _GEN_4123; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4322 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ftq_idx : _GEN_4124; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4323 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_br_tag : _GEN_4125; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4324 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_br_mask : _GEN_4126; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4325 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_sfb : _GEN_4127; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4326 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_jal : _GEN_4128; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4327 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_jalr : _GEN_4129; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4328 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_br : _GEN_4130; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4329 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_iw_p2_poisoned : _GEN_4131; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4330 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_iw_p1_poisoned : _GEN_4132; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4331 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_iw_state : _GEN_4133; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4332 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_op3_sel : _GEN_4134; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4333 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_is_std : _GEN_4135; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4334 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_is_sta : _GEN_4136; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4335 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_is_load : _GEN_4137; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4336 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_csr_cmd : _GEN_4138; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4337 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_fcn_dw : _GEN_4139; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4338 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_op_fcn : _GEN_4140; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4339 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_imm_sel : _GEN_4141; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4340 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_op2_sel : _GEN_4142; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4341 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_op1_sel : _GEN_4143; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4342 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_ctrl_br_type : _GEN_4144; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4343 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_fu_code : _GEN_4145; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4344 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_iq_type : _GEN_4146; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_4345 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_debug_pc : _GEN_4147; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4346 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_rvc : _GEN_4148; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4347 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_debug_inst : _GEN_4149; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4348 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_inst : _GEN_4150; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4349 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_uopc : _GEN_4151; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4350 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_address_num : _GEN_4152; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4351 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_rob_inst_idx : _GEN_4153; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4352 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_self_index : _GEN_4154; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4353 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_split_num : _GEN_4155; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4354 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_op2_sel : _GEN_4156; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4355 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_op1_sel : _GEN_4157; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4356 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_stale_pflag : _GEN_4158; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4357 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_pflag_busy : _GEN_4159; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4358 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_pwflag : _GEN_4160; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4359 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_prflag : _GEN_4161; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4360 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_wflag : _GEN_4162; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4361 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_rflag : _GEN_4163; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4362 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_lrs3_rtype : _GEN_4164; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4363 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_shift : _GEN_4165; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4364 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_is_unicore : _GEN_4166; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4365 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_switch_off : _GEN_4167; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4366 = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) ?
    issue_slots_1_uop_switch : _GEN_4168; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_debug_tsrc = slots_2_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4369 = _T_485 ? issue_slots_2_uop_debug_tsrc : _GEN_4171; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_debug_fsrc = slots_2_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4370 = _T_485 ? issue_slots_2_uop_debug_fsrc : _GEN_4172; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_bp_xcpt_if = slots_2_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4371 = _T_485 ? issue_slots_2_uop_bp_xcpt_if : _GEN_4173; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_bp_debug_if = slots_2_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4372 = _T_485 ? issue_slots_2_uop_bp_debug_if : _GEN_4174; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_xcpt_ma_if = slots_2_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4373 = _T_485 ? issue_slots_2_uop_xcpt_ma_if : _GEN_4175; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_xcpt_ae_if = slots_2_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4374 = _T_485 ? issue_slots_2_uop_xcpt_ae_if : _GEN_4176; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_xcpt_pf_if = slots_2_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4375 = _T_485 ? issue_slots_2_uop_xcpt_pf_if : _GEN_4177; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_fp_single = slots_2_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4376 = _T_485 ? issue_slots_2_uop_fp_single : _GEN_4178; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_fp_val = slots_2_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4377 = _T_485 ? issue_slots_2_uop_fp_val : _GEN_4179; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_frs3_en = slots_2_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4378 = _T_485 ? issue_slots_2_uop_frs3_en : _GEN_4180; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_lrs2_rtype = slots_2_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4379 = _T_485 ? issue_slots_2_uop_lrs2_rtype : _GEN_4181; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_lrs1_rtype = slots_2_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4380 = _T_485 ? issue_slots_2_uop_lrs1_rtype : _GEN_4182; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_dst_rtype = slots_2_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4381 = _T_485 ? issue_slots_2_uop_dst_rtype : _GEN_4183; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ldst_val = slots_2_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4382 = _T_485 ? issue_slots_2_uop_ldst_val : _GEN_4184; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_lrs3 = slots_2_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4383 = _T_485 ? issue_slots_2_uop_lrs3 : _GEN_4185; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_lrs2 = slots_2_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4384 = _T_485 ? issue_slots_2_uop_lrs2 : _GEN_4186; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_lrs1 = slots_2_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4385 = _T_485 ? issue_slots_2_uop_lrs1 : _GEN_4187; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_ldst = slots_2_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4386 = _T_485 ? issue_slots_2_uop_ldst : _GEN_4188; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ldst_is_rs1 = slots_2_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4387 = _T_485 ? issue_slots_2_uop_ldst_is_rs1 : _GEN_4189; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_flush_on_commit = slots_2_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4388 = _T_485 ? issue_slots_2_uop_flush_on_commit : _GEN_4190; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_unique = slots_2_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4389 = _T_485 ? issue_slots_2_uop_is_unique : _GEN_4191; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_sys_pc2epc = slots_2_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4390 = _T_485 ? issue_slots_2_uop_is_sys_pc2epc : _GEN_4192; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_uses_stq = slots_2_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4391 = _T_485 ? issue_slots_2_uop_uses_stq : _GEN_4193; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_uses_ldq = slots_2_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4392 = _T_485 ? issue_slots_2_uop_uses_ldq : _GEN_4194; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_amo = slots_2_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4393 = _T_485 ? issue_slots_2_uop_is_amo : _GEN_4195; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_fencei = slots_2_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4394 = _T_485 ? issue_slots_2_uop_is_fencei : _GEN_4196; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_fence = slots_2_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4395 = _T_485 ? issue_slots_2_uop_is_fence : _GEN_4197; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_mem_signed = slots_2_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4396 = _T_485 ? issue_slots_2_uop_mem_signed : _GEN_4198; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_mem_size = slots_2_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4397 = _T_485 ? issue_slots_2_uop_mem_size : _GEN_4199; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_mem_cmd = slots_2_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4398 = _T_485 ? issue_slots_2_uop_mem_cmd : _GEN_4200; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_bypassable = slots_2_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4399 = _T_485 ? issue_slots_2_uop_bypassable : _GEN_4201; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_2_uop_exc_cause = slots_2_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4400 = _T_485 ? issue_slots_2_uop_exc_cause : _GEN_4202; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_exception = slots_2_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4401 = _T_485 ? issue_slots_2_uop_exception : _GEN_4203; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_stale_pdst = slots_2_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4402 = _T_485 ? issue_slots_2_uop_stale_pdst : _GEN_4204; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ppred_busy = slots_2_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4403 = _T_485 ? issue_slots_2_uop_ppred_busy : _GEN_4205; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_prs3_busy = slots_2_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4404 = _T_485 ? issue_slots_2_uop_prs3_busy : _GEN_4206; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_prs2_busy = slots_2_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4405 = _T_485 ? issue_slots_2_uop_prs2_busy : _GEN_4207; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_prs1_busy = slots_2_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4406 = _T_485 ? issue_slots_2_uop_prs1_busy : _GEN_4208; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_ppred = slots_2_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4407 = _T_485 ? issue_slots_2_uop_ppred : _GEN_4209; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_prs3 = slots_2_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4408 = _T_485 ? issue_slots_2_uop_prs3 : _GEN_4210; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_prs2 = slots_2_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4409 = _T_485 ? issue_slots_2_uop_prs2 : _GEN_4211; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_prs1 = slots_2_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4410 = _T_485 ? issue_slots_2_uop_prs1 : _GEN_4212; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_pdst = slots_2_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4411 = _T_485 ? issue_slots_2_uop_pdst : _GEN_4213; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_rxq_idx = slots_2_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4412 = _T_485 ? issue_slots_2_uop_rxq_idx : _GEN_4214; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_stq_idx = slots_2_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4413 = _T_485 ? issue_slots_2_uop_stq_idx : _GEN_4215; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_ldq_idx = slots_2_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4414 = _T_485 ? issue_slots_2_uop_ldq_idx : _GEN_4216; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_rob_idx = slots_2_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4415 = _T_485 ? issue_slots_2_uop_rob_idx : _GEN_4217; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_2_uop_csr_addr = slots_2_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4416 = _T_485 ? issue_slots_2_uop_csr_addr : _GEN_4218; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_2_uop_imm_packed = slots_2_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4417 = _T_485 ? issue_slots_2_uop_imm_packed : _GEN_4219; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_taken = slots_2_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4418 = _T_485 ? issue_slots_2_uop_taken : _GEN_4220; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_pc_lob = slots_2_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4419 = _T_485 ? issue_slots_2_uop_pc_lob : _GEN_4221; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_edge_inst = slots_2_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4420 = _T_485 ? issue_slots_2_uop_edge_inst : _GEN_4222; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_ftq_idx = slots_2_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4421 = _T_485 ? issue_slots_2_uop_ftq_idx : _GEN_4223; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_br_tag = slots_2_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4422 = _T_485 ? issue_slots_2_uop_br_tag : _GEN_4224; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_2_uop_br_mask = slots_2_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4423 = _T_485 ? issue_slots_2_uop_br_mask : _GEN_4225; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_sfb = slots_2_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4424 = _T_485 ? issue_slots_2_uop_is_sfb : _GEN_4226; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_jal = slots_2_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4425 = _T_485 ? issue_slots_2_uop_is_jal : _GEN_4227; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_jalr = slots_2_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4426 = _T_485 ? issue_slots_2_uop_is_jalr : _GEN_4228; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_br = slots_2_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4427 = _T_485 ? issue_slots_2_uop_is_br : _GEN_4229; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_iw_p2_poisoned = slots_2_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4428 = _T_485 ? issue_slots_2_uop_iw_p2_poisoned : _GEN_4230; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_iw_p1_poisoned = slots_2_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4429 = _T_485 ? issue_slots_2_uop_iw_p1_poisoned : _GEN_4231; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_iw_state = slots_2_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4430 = _T_485 ? issue_slots_2_uop_iw_state : _GEN_4232; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_ctrl_op3_sel = slots_2_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4431 = _T_485 ? issue_slots_2_uop_ctrl_op3_sel : _GEN_4233; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_is_std = slots_2_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4432 = _T_485 ? issue_slots_2_uop_ctrl_is_std : _GEN_4234; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_is_sta = slots_2_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4433 = _T_485 ? issue_slots_2_uop_ctrl_is_sta : _GEN_4235; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_is_load = slots_2_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4434 = _T_485 ? issue_slots_2_uop_ctrl_is_load : _GEN_4236; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_ctrl_csr_cmd = slots_2_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4435 = _T_485 ? issue_slots_2_uop_ctrl_csr_cmd : _GEN_4237; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_fcn_dw = slots_2_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4436 = _T_485 ? issue_slots_2_uop_ctrl_fcn_dw : _GEN_4238; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_ctrl_op_fcn = slots_2_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4437 = _T_485 ? issue_slots_2_uop_ctrl_op_fcn : _GEN_4239; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_ctrl_imm_sel = slots_2_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4438 = _T_485 ? issue_slots_2_uop_ctrl_imm_sel : _GEN_4240; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_ctrl_op2_sel = slots_2_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4439 = _T_485 ? issue_slots_2_uop_ctrl_op2_sel : _GEN_4241; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_ctrl_op1_sel = slots_2_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4440 = _T_485 ? issue_slots_2_uop_ctrl_op1_sel : _GEN_4242; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_ctrl_br_type = slots_2_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4441 = _T_485 ? issue_slots_2_uop_ctrl_br_type : _GEN_4243; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4442 = _T_485 ? issue_slots_2_uop_fu_code : _GEN_4244; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_iq_type = slots_2_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4443 = _T_485 ? issue_slots_2_uop_iq_type : _GEN_4245; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_2_uop_debug_pc = slots_2_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4444 = _T_485 ? issue_slots_2_uop_debug_pc : _GEN_4246; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_rvc = slots_2_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4445 = _T_485 ? issue_slots_2_uop_is_rvc : _GEN_4247; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_2_uop_debug_inst = slots_2_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4446 = _T_485 ? issue_slots_2_uop_debug_inst : _GEN_4248; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_2_uop_inst = slots_2_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4447 = _T_485 ? issue_slots_2_uop_inst : _GEN_4249; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_uopc = slots_2_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4448 = _T_485 ? issue_slots_2_uop_uopc : _GEN_4250; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_address_num = slots_2_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4449 = _T_485 ? issue_slots_2_uop_address_num : _GEN_4251; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_rob_inst_idx = slots_2_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4450 = _T_485 ? issue_slots_2_uop_rob_inst_idx : _GEN_4252; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_self_index = slots_2_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4451 = _T_485 ? issue_slots_2_uop_self_index : _GEN_4253; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_split_num = slots_2_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4452 = _T_485 ? issue_slots_2_uop_split_num : _GEN_4254; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_op2_sel = slots_2_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4453 = _T_485 ? issue_slots_2_uop_op2_sel : _GEN_4255; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_op1_sel = slots_2_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4454 = _T_485 ? issue_slots_2_uop_op1_sel : _GEN_4256; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_stale_pflag = slots_2_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4455 = _T_485 ? issue_slots_2_uop_stale_pflag : _GEN_4257; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_pflag_busy = slots_2_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4456 = _T_485 ? issue_slots_2_uop_pflag_busy : _GEN_4258; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_pwflag = slots_2_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4457 = _T_485 ? issue_slots_2_uop_pwflag : _GEN_4259; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_prflag = slots_2_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4458 = _T_485 ? issue_slots_2_uop_prflag : _GEN_4260; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_wflag = slots_2_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4459 = _T_485 ? issue_slots_2_uop_wflag : _GEN_4261; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_rflag = slots_2_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4460 = _T_485 ? issue_slots_2_uop_rflag : _GEN_4262; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_lrs3_rtype = slots_2_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4461 = _T_485 ? issue_slots_2_uop_lrs3_rtype : _GEN_4263; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_shift = slots_2_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4462 = _T_485 ? issue_slots_2_uop_shift : _GEN_4264; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_unicore = slots_2_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4463 = _T_485 ? issue_slots_2_uop_is_unicore : _GEN_4265; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_switch_off = slots_2_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4464 = _T_485 ? issue_slots_2_uop_switch_off : _GEN_4266; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_switch = slots_2_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4465 = _T_485 ? issue_slots_2_uop_switch : _GEN_4267; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4468 = _T_496 & ~_T_467 ? issue_slots_2_uop_debug_tsrc : _GEN_4270; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4469 = _T_496 & ~_T_467 ? issue_slots_2_uop_debug_fsrc : _GEN_4271; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4470 = _T_496 & ~_T_467 ? issue_slots_2_uop_bp_xcpt_if : _GEN_4272; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4471 = _T_496 & ~_T_467 ? issue_slots_2_uop_bp_debug_if : _GEN_4273; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4472 = _T_496 & ~_T_467 ? issue_slots_2_uop_xcpt_ma_if : _GEN_4274; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4473 = _T_496 & ~_T_467 ? issue_slots_2_uop_xcpt_ae_if : _GEN_4275; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4474 = _T_496 & ~_T_467 ? issue_slots_2_uop_xcpt_pf_if : _GEN_4276; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4475 = _T_496 & ~_T_467 ? issue_slots_2_uop_fp_single : _GEN_4277; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4476 = _T_496 & ~_T_467 ? issue_slots_2_uop_fp_val : _GEN_4278; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4477 = _T_496 & ~_T_467 ? issue_slots_2_uop_frs3_en : _GEN_4279; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4478 = _T_496 & ~_T_467 ? issue_slots_2_uop_lrs2_rtype : _GEN_4280; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4479 = _T_496 & ~_T_467 ? issue_slots_2_uop_lrs1_rtype : _GEN_4281; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4480 = _T_496 & ~_T_467 ? issue_slots_2_uop_dst_rtype : _GEN_4282; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4481 = _T_496 & ~_T_467 ? issue_slots_2_uop_ldst_val : _GEN_4283; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4482 = _T_496 & ~_T_467 ? issue_slots_2_uop_lrs3 : _GEN_4284; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4483 = _T_496 & ~_T_467 ? issue_slots_2_uop_lrs2 : _GEN_4285; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4484 = _T_496 & ~_T_467 ? issue_slots_2_uop_lrs1 : _GEN_4286; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4485 = _T_496 & ~_T_467 ? issue_slots_2_uop_ldst : _GEN_4287; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4486 = _T_496 & ~_T_467 ? issue_slots_2_uop_ldst_is_rs1 : _GEN_4288; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4487 = _T_496 & ~_T_467 ? issue_slots_2_uop_flush_on_commit : _GEN_4289; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4488 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_unique : _GEN_4290; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4489 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_sys_pc2epc : _GEN_4291; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4490 = _T_496 & ~_T_467 ? issue_slots_2_uop_uses_stq : _GEN_4292; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4491 = _T_496 & ~_T_467 ? issue_slots_2_uop_uses_ldq : _GEN_4293; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4492 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_amo : _GEN_4294; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4493 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_fencei : _GEN_4295; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4494 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_fence : _GEN_4296; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4495 = _T_496 & ~_T_467 ? issue_slots_2_uop_mem_signed : _GEN_4297; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4496 = _T_496 & ~_T_467 ? issue_slots_2_uop_mem_size : _GEN_4298; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4497 = _T_496 & ~_T_467 ? issue_slots_2_uop_mem_cmd : _GEN_4299; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4498 = _T_496 & ~_T_467 ? issue_slots_2_uop_bypassable : _GEN_4300; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_4499 = _T_496 & ~_T_467 ? issue_slots_2_uop_exc_cause : _GEN_4301; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4500 = _T_496 & ~_T_467 ? issue_slots_2_uop_exception : _GEN_4302; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4501 = _T_496 & ~_T_467 ? issue_slots_2_uop_stale_pdst : _GEN_4303; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4502 = _T_496 & ~_T_467 ? issue_slots_2_uop_ppred_busy : _GEN_4304; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4503 = _T_496 & ~_T_467 ? issue_slots_2_uop_prs3_busy : _GEN_4305; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4504 = _T_496 & ~_T_467 ? issue_slots_2_uop_prs2_busy : _GEN_4306; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4505 = _T_496 & ~_T_467 ? issue_slots_2_uop_prs1_busy : _GEN_4307; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4506 = _T_496 & ~_T_467 ? issue_slots_2_uop_ppred : _GEN_4308; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4507 = _T_496 & ~_T_467 ? issue_slots_2_uop_prs3 : _GEN_4309; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4508 = _T_496 & ~_T_467 ? issue_slots_2_uop_prs2 : _GEN_4310; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4509 = _T_496 & ~_T_467 ? issue_slots_2_uop_prs1 : _GEN_4311; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4510 = _T_496 & ~_T_467 ? issue_slots_2_uop_pdst : _GEN_4312; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4511 = _T_496 & ~_T_467 ? issue_slots_2_uop_rxq_idx : _GEN_4313; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4512 = _T_496 & ~_T_467 ? issue_slots_2_uop_stq_idx : _GEN_4314; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4513 = _T_496 & ~_T_467 ? issue_slots_2_uop_ldq_idx : _GEN_4315; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4514 = _T_496 & ~_T_467 ? issue_slots_2_uop_rob_idx : _GEN_4316; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4515 = _T_496 & ~_T_467 ? issue_slots_2_uop_csr_addr : _GEN_4317; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_4516 = _T_496 & ~_T_467 ? issue_slots_2_uop_imm_packed : _GEN_4318; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4517 = _T_496 & ~_T_467 ? issue_slots_2_uop_taken : _GEN_4319; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4518 = _T_496 & ~_T_467 ? issue_slots_2_uop_pc_lob : _GEN_4320; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4519 = _T_496 & ~_T_467 ? issue_slots_2_uop_edge_inst : _GEN_4321; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4520 = _T_496 & ~_T_467 ? issue_slots_2_uop_ftq_idx : _GEN_4322; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4521 = _T_496 & ~_T_467 ? issue_slots_2_uop_br_tag : _GEN_4323; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4522 = _T_496 & ~_T_467 ? issue_slots_2_uop_br_mask : _GEN_4324; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4523 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_sfb : _GEN_4325; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4524 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_jal : _GEN_4326; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4525 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_jalr : _GEN_4327; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4526 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_br : _GEN_4328; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4527 = _T_496 & ~_T_467 ? issue_slots_2_uop_iw_p2_poisoned : _GEN_4329; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4528 = _T_496 & ~_T_467 ? issue_slots_2_uop_iw_p1_poisoned : _GEN_4330; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4529 = _T_496 & ~_T_467 ? issue_slots_2_uop_iw_state : _GEN_4331; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4530 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_op3_sel : _GEN_4332; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4531 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_is_std : _GEN_4333; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4532 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_is_sta : _GEN_4334; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4533 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_is_load : _GEN_4335; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4534 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_csr_cmd : _GEN_4336; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4535 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_fcn_dw : _GEN_4337; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4536 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_op_fcn : _GEN_4338; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4537 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_imm_sel : _GEN_4339; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4538 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_op2_sel : _GEN_4340; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4539 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_op1_sel : _GEN_4341; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4540 = _T_496 & ~_T_467 ? issue_slots_2_uop_ctrl_br_type : _GEN_4342; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4541 = _T_496 & ~_T_467 ? issue_slots_2_uop_fu_code : _GEN_4343; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4542 = _T_496 & ~_T_467 ? issue_slots_2_uop_iq_type : _GEN_4344; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_4543 = _T_496 & ~_T_467 ? issue_slots_2_uop_debug_pc : _GEN_4345; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4544 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_rvc : _GEN_4346; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4545 = _T_496 & ~_T_467 ? issue_slots_2_uop_debug_inst : _GEN_4347; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4546 = _T_496 & ~_T_467 ? issue_slots_2_uop_inst : _GEN_4348; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4547 = _T_496 & ~_T_467 ? issue_slots_2_uop_uopc : _GEN_4349; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4548 = _T_496 & ~_T_467 ? issue_slots_2_uop_address_num : _GEN_4350; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4549 = _T_496 & ~_T_467 ? issue_slots_2_uop_rob_inst_idx : _GEN_4351; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4550 = _T_496 & ~_T_467 ? issue_slots_2_uop_self_index : _GEN_4352; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4551 = _T_496 & ~_T_467 ? issue_slots_2_uop_split_num : _GEN_4353; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4552 = _T_496 & ~_T_467 ? issue_slots_2_uop_op2_sel : _GEN_4354; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4553 = _T_496 & ~_T_467 ? issue_slots_2_uop_op1_sel : _GEN_4355; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4554 = _T_496 & ~_T_467 ? issue_slots_2_uop_stale_pflag : _GEN_4356; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4555 = _T_496 & ~_T_467 ? issue_slots_2_uop_pflag_busy : _GEN_4357; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4556 = _T_496 & ~_T_467 ? issue_slots_2_uop_pwflag : _GEN_4358; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4557 = _T_496 & ~_T_467 ? issue_slots_2_uop_prflag : _GEN_4359; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4558 = _T_496 & ~_T_467 ? issue_slots_2_uop_wflag : _GEN_4360; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4559 = _T_496 & ~_T_467 ? issue_slots_2_uop_rflag : _GEN_4361; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4560 = _T_496 & ~_T_467 ? issue_slots_2_uop_lrs3_rtype : _GEN_4362; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4561 = _T_496 & ~_T_467 ? issue_slots_2_uop_shift : _GEN_4363; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4562 = _T_496 & ~_T_467 ? issue_slots_2_uop_is_unicore : _GEN_4364; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4563 = _T_496 & ~_T_467 ? issue_slots_2_uop_switch_off : _GEN_4365; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4564 = _T_496 & ~_T_467 ? issue_slots_2_uop_switch : _GEN_4366; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_debug_tsrc = slots_3_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4567 = _T_515 ? issue_slots_3_uop_debug_tsrc : _GEN_4369; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_debug_fsrc = slots_3_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4568 = _T_515 ? issue_slots_3_uop_debug_fsrc : _GEN_4370; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_bp_xcpt_if = slots_3_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4569 = _T_515 ? issue_slots_3_uop_bp_xcpt_if : _GEN_4371; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_bp_debug_if = slots_3_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4570 = _T_515 ? issue_slots_3_uop_bp_debug_if : _GEN_4372; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_xcpt_ma_if = slots_3_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4571 = _T_515 ? issue_slots_3_uop_xcpt_ma_if : _GEN_4373; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_xcpt_ae_if = slots_3_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4572 = _T_515 ? issue_slots_3_uop_xcpt_ae_if : _GEN_4374; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_xcpt_pf_if = slots_3_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4573 = _T_515 ? issue_slots_3_uop_xcpt_pf_if : _GEN_4375; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_fp_single = slots_3_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4574 = _T_515 ? issue_slots_3_uop_fp_single : _GEN_4376; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_fp_val = slots_3_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4575 = _T_515 ? issue_slots_3_uop_fp_val : _GEN_4377; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_frs3_en = slots_3_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4576 = _T_515 ? issue_slots_3_uop_frs3_en : _GEN_4378; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_lrs2_rtype = slots_3_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4577 = _T_515 ? issue_slots_3_uop_lrs2_rtype : _GEN_4379; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_lrs1_rtype = slots_3_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4578 = _T_515 ? issue_slots_3_uop_lrs1_rtype : _GEN_4380; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_dst_rtype = slots_3_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4579 = _T_515 ? issue_slots_3_uop_dst_rtype : _GEN_4381; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ldst_val = slots_3_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4580 = _T_515 ? issue_slots_3_uop_ldst_val : _GEN_4382; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_lrs3 = slots_3_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4581 = _T_515 ? issue_slots_3_uop_lrs3 : _GEN_4383; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_lrs2 = slots_3_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4582 = _T_515 ? issue_slots_3_uop_lrs2 : _GEN_4384; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_lrs1 = slots_3_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4583 = _T_515 ? issue_slots_3_uop_lrs1 : _GEN_4385; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_ldst = slots_3_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4584 = _T_515 ? issue_slots_3_uop_ldst : _GEN_4386; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ldst_is_rs1 = slots_3_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4585 = _T_515 ? issue_slots_3_uop_ldst_is_rs1 : _GEN_4387; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_flush_on_commit = slots_3_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4586 = _T_515 ? issue_slots_3_uop_flush_on_commit : _GEN_4388; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_unique = slots_3_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4587 = _T_515 ? issue_slots_3_uop_is_unique : _GEN_4389; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_sys_pc2epc = slots_3_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4588 = _T_515 ? issue_slots_3_uop_is_sys_pc2epc : _GEN_4390; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_uses_stq = slots_3_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4589 = _T_515 ? issue_slots_3_uop_uses_stq : _GEN_4391; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_uses_ldq = slots_3_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4590 = _T_515 ? issue_slots_3_uop_uses_ldq : _GEN_4392; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_amo = slots_3_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4591 = _T_515 ? issue_slots_3_uop_is_amo : _GEN_4393; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_fencei = slots_3_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4592 = _T_515 ? issue_slots_3_uop_is_fencei : _GEN_4394; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_fence = slots_3_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4593 = _T_515 ? issue_slots_3_uop_is_fence : _GEN_4395; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_mem_signed = slots_3_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4594 = _T_515 ? issue_slots_3_uop_mem_signed : _GEN_4396; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_mem_size = slots_3_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4595 = _T_515 ? issue_slots_3_uop_mem_size : _GEN_4397; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_mem_cmd = slots_3_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4596 = _T_515 ? issue_slots_3_uop_mem_cmd : _GEN_4398; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_bypassable = slots_3_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4597 = _T_515 ? issue_slots_3_uop_bypassable : _GEN_4399; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_3_uop_exc_cause = slots_3_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4598 = _T_515 ? issue_slots_3_uop_exc_cause : _GEN_4400; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_exception = slots_3_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4599 = _T_515 ? issue_slots_3_uop_exception : _GEN_4401; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_stale_pdst = slots_3_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4600 = _T_515 ? issue_slots_3_uop_stale_pdst : _GEN_4402; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ppred_busy = slots_3_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4601 = _T_515 ? issue_slots_3_uop_ppred_busy : _GEN_4403; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_prs3_busy = slots_3_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4602 = _T_515 ? issue_slots_3_uop_prs3_busy : _GEN_4404; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_prs2_busy = slots_3_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4603 = _T_515 ? issue_slots_3_uop_prs2_busy : _GEN_4405; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_prs1_busy = slots_3_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4604 = _T_515 ? issue_slots_3_uop_prs1_busy : _GEN_4406; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_ppred = slots_3_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4605 = _T_515 ? issue_slots_3_uop_ppred : _GEN_4407; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_prs3 = slots_3_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4606 = _T_515 ? issue_slots_3_uop_prs3 : _GEN_4408; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_prs2 = slots_3_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4607 = _T_515 ? issue_slots_3_uop_prs2 : _GEN_4409; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_prs1 = slots_3_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4608 = _T_515 ? issue_slots_3_uop_prs1 : _GEN_4410; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_pdst = slots_3_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4609 = _T_515 ? issue_slots_3_uop_pdst : _GEN_4411; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_rxq_idx = slots_3_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4610 = _T_515 ? issue_slots_3_uop_rxq_idx : _GEN_4412; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_stq_idx = slots_3_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4611 = _T_515 ? issue_slots_3_uop_stq_idx : _GEN_4413; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_ldq_idx = slots_3_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4612 = _T_515 ? issue_slots_3_uop_ldq_idx : _GEN_4414; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_rob_idx = slots_3_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4613 = _T_515 ? issue_slots_3_uop_rob_idx : _GEN_4415; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_3_uop_csr_addr = slots_3_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4614 = _T_515 ? issue_slots_3_uop_csr_addr : _GEN_4416; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_3_uop_imm_packed = slots_3_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4615 = _T_515 ? issue_slots_3_uop_imm_packed : _GEN_4417; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_taken = slots_3_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4616 = _T_515 ? issue_slots_3_uop_taken : _GEN_4418; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_pc_lob = slots_3_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4617 = _T_515 ? issue_slots_3_uop_pc_lob : _GEN_4419; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_edge_inst = slots_3_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4618 = _T_515 ? issue_slots_3_uop_edge_inst : _GEN_4420; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_ftq_idx = slots_3_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4619 = _T_515 ? issue_slots_3_uop_ftq_idx : _GEN_4421; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_br_tag = slots_3_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4620 = _T_515 ? issue_slots_3_uop_br_tag : _GEN_4422; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_3_uop_br_mask = slots_3_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4621 = _T_515 ? issue_slots_3_uop_br_mask : _GEN_4423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_sfb = slots_3_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4622 = _T_515 ? issue_slots_3_uop_is_sfb : _GEN_4424; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_jal = slots_3_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4623 = _T_515 ? issue_slots_3_uop_is_jal : _GEN_4425; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_jalr = slots_3_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4624 = _T_515 ? issue_slots_3_uop_is_jalr : _GEN_4426; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_br = slots_3_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4625 = _T_515 ? issue_slots_3_uop_is_br : _GEN_4427; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_iw_p2_poisoned = slots_3_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4626 = _T_515 ? issue_slots_3_uop_iw_p2_poisoned : _GEN_4428; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_iw_p1_poisoned = slots_3_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4627 = _T_515 ? issue_slots_3_uop_iw_p1_poisoned : _GEN_4429; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_iw_state = slots_3_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4628 = _T_515 ? issue_slots_3_uop_iw_state : _GEN_4430; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_ctrl_op3_sel = slots_3_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4629 = _T_515 ? issue_slots_3_uop_ctrl_op3_sel : _GEN_4431; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_is_std = slots_3_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4630 = _T_515 ? issue_slots_3_uop_ctrl_is_std : _GEN_4432; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_is_sta = slots_3_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4631 = _T_515 ? issue_slots_3_uop_ctrl_is_sta : _GEN_4433; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_is_load = slots_3_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4632 = _T_515 ? issue_slots_3_uop_ctrl_is_load : _GEN_4434; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_ctrl_csr_cmd = slots_3_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4633 = _T_515 ? issue_slots_3_uop_ctrl_csr_cmd : _GEN_4435; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_fcn_dw = slots_3_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4634 = _T_515 ? issue_slots_3_uop_ctrl_fcn_dw : _GEN_4436; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_ctrl_op_fcn = slots_3_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4635 = _T_515 ? issue_slots_3_uop_ctrl_op_fcn : _GEN_4437; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_ctrl_imm_sel = slots_3_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4636 = _T_515 ? issue_slots_3_uop_ctrl_imm_sel : _GEN_4438; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_ctrl_op2_sel = slots_3_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4637 = _T_515 ? issue_slots_3_uop_ctrl_op2_sel : _GEN_4439; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_ctrl_op1_sel = slots_3_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4638 = _T_515 ? issue_slots_3_uop_ctrl_op1_sel : _GEN_4440; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_ctrl_br_type = slots_3_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4639 = _T_515 ? issue_slots_3_uop_ctrl_br_type : _GEN_4441; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4640 = _T_515 ? issue_slots_3_uop_fu_code : _GEN_4442; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_iq_type = slots_3_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4641 = _T_515 ? issue_slots_3_uop_iq_type : _GEN_4443; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_3_uop_debug_pc = slots_3_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4642 = _T_515 ? issue_slots_3_uop_debug_pc : _GEN_4444; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_rvc = slots_3_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4643 = _T_515 ? issue_slots_3_uop_is_rvc : _GEN_4445; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_3_uop_debug_inst = slots_3_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4644 = _T_515 ? issue_slots_3_uop_debug_inst : _GEN_4446; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_3_uop_inst = slots_3_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4645 = _T_515 ? issue_slots_3_uop_inst : _GEN_4447; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_uopc = slots_3_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4646 = _T_515 ? issue_slots_3_uop_uopc : _GEN_4448; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_address_num = slots_3_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4647 = _T_515 ? issue_slots_3_uop_address_num : _GEN_4449; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_rob_inst_idx = slots_3_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4648 = _T_515 ? issue_slots_3_uop_rob_inst_idx : _GEN_4450; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_self_index = slots_3_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4649 = _T_515 ? issue_slots_3_uop_self_index : _GEN_4451; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_split_num = slots_3_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4650 = _T_515 ? issue_slots_3_uop_split_num : _GEN_4452; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_op2_sel = slots_3_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4651 = _T_515 ? issue_slots_3_uop_op2_sel : _GEN_4453; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_op1_sel = slots_3_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4652 = _T_515 ? issue_slots_3_uop_op1_sel : _GEN_4454; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_stale_pflag = slots_3_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4653 = _T_515 ? issue_slots_3_uop_stale_pflag : _GEN_4455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_pflag_busy = slots_3_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4654 = _T_515 ? issue_slots_3_uop_pflag_busy : _GEN_4456; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_pwflag = slots_3_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4655 = _T_515 ? issue_slots_3_uop_pwflag : _GEN_4457; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_prflag = slots_3_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4656 = _T_515 ? issue_slots_3_uop_prflag : _GEN_4458; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_wflag = slots_3_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4657 = _T_515 ? issue_slots_3_uop_wflag : _GEN_4459; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_rflag = slots_3_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4658 = _T_515 ? issue_slots_3_uop_rflag : _GEN_4460; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_lrs3_rtype = slots_3_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4659 = _T_515 ? issue_slots_3_uop_lrs3_rtype : _GEN_4461; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_shift = slots_3_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4660 = _T_515 ? issue_slots_3_uop_shift : _GEN_4462; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_unicore = slots_3_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4661 = _T_515 ? issue_slots_3_uop_is_unicore : _GEN_4463; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_switch_off = slots_3_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4662 = _T_515 ? issue_slots_3_uop_switch_off : _GEN_4464; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_switch = slots_3_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4663 = _T_515 ? issue_slots_3_uop_switch : _GEN_4465; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4666 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_debug_tsrc : _GEN_4468; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4667 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_debug_fsrc : _GEN_4469; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4668 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_bp_xcpt_if : _GEN_4470; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4669 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_bp_debug_if : _GEN_4471; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4670 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_xcpt_ma_if : _GEN_4472; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4671 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_xcpt_ae_if : _GEN_4473; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4672 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_xcpt_pf_if : _GEN_4474; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4673 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_fp_single : _GEN_4475; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4674 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_fp_val : _GEN_4476; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4675 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_frs3_en : _GEN_4477; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4676 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_lrs2_rtype : _GEN_4478; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4677 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_lrs1_rtype : _GEN_4479; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4678 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_dst_rtype : _GEN_4480; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4679 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ldst_val : _GEN_4481; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4680 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_lrs3 : _GEN_4482; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4681 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_lrs2 : _GEN_4483; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4682 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_lrs1 : _GEN_4484; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4683 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ldst : _GEN_4485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4684 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ldst_is_rs1 : _GEN_4486; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4685 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_flush_on_commit : _GEN_4487; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4686 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_unique : _GEN_4488; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4687 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_sys_pc2epc : _GEN_4489; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4688 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_uses_stq : _GEN_4490; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4689 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_uses_ldq : _GEN_4491; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4690 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_amo : _GEN_4492; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4691 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_fencei : _GEN_4493; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4692 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_fence : _GEN_4494; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4693 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_mem_signed : _GEN_4495; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4694 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_mem_size : _GEN_4496; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4695 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_mem_cmd : _GEN_4497; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4696 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_bypassable : _GEN_4498; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_4697 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_exc_cause : _GEN_4499; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4698 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_exception : _GEN_4500; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4699 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_stale_pdst : _GEN_4501; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4700 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ppred_busy : _GEN_4502; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4701 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_prs3_busy : _GEN_4503; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4702 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_prs2_busy : _GEN_4504; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4703 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_prs1_busy : _GEN_4505; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4704 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ppred : _GEN_4506; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4705 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_prs3 : _GEN_4507; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4706 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_prs2 : _GEN_4508; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4707 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_prs1 : _GEN_4509; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4708 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_pdst : _GEN_4510; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4709 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_rxq_idx : _GEN_4511; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4710 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_stq_idx : _GEN_4512; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4711 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ldq_idx : _GEN_4513; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4712 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_rob_idx : _GEN_4514; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4713 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_csr_addr : _GEN_4515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_4714 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_imm_packed : _GEN_4516; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4715 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_taken : _GEN_4517; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4716 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_pc_lob : _GEN_4518; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4717 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_edge_inst : _GEN_4519; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4718 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ftq_idx : _GEN_4520; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4719 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_br_tag : _GEN_4521; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4720 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_br_mask : _GEN_4522; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4721 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_sfb : _GEN_4523; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4722 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_jal : _GEN_4524; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4723 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_jalr : _GEN_4525; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4724 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_br : _GEN_4526; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4725 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_iw_p2_poisoned : _GEN_4527; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4726 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_iw_p1_poisoned : _GEN_4528; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4727 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_iw_state : _GEN_4529; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4728 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_op3_sel : _GEN_4530
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4729 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_is_std : _GEN_4531; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4730 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_is_sta : _GEN_4532; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4731 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_is_load : _GEN_4533; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4732 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_csr_cmd : _GEN_4534
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4733 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_fcn_dw : _GEN_4535; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4734 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_op_fcn : _GEN_4536; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4735 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_imm_sel : _GEN_4537
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4736 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_op2_sel : _GEN_4538
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4737 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_op1_sel : _GEN_4539
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4738 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_ctrl_br_type : _GEN_4540
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4739 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_fu_code : _GEN_4541; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4740 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_iq_type : _GEN_4542; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_4741 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_debug_pc : _GEN_4543; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4742 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_rvc : _GEN_4544; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4743 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_debug_inst : _GEN_4545; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4744 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_inst : _GEN_4546; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4745 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_uopc : _GEN_4547; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4746 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_address_num : _GEN_4548; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4747 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_rob_inst_idx : _GEN_4549
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4748 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_self_index : _GEN_4550; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4749 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_split_num : _GEN_4551; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4750 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_op2_sel : _GEN_4552; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4751 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_op1_sel : _GEN_4553; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4752 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_stale_pflag : _GEN_4554; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4753 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_pflag_busy : _GEN_4555; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4754 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_pwflag : _GEN_4556; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4755 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_prflag : _GEN_4557; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4756 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_wflag : _GEN_4558; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4757 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_rflag : _GEN_4559; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4758 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_lrs3_rtype : _GEN_4560; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4759 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_shift : _GEN_4561; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4760 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_is_unicore : _GEN_4562; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4761 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_switch_off : _GEN_4563; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4762 = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 ? issue_slots_3_uop_switch : _GEN_4564; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_debug_tsrc = slots_4_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4765 = _T_545 ? issue_slots_4_uop_debug_tsrc : _GEN_4567; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_debug_fsrc = slots_4_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4766 = _T_545 ? issue_slots_4_uop_debug_fsrc : _GEN_4568; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_bp_xcpt_if = slots_4_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4767 = _T_545 ? issue_slots_4_uop_bp_xcpt_if : _GEN_4569; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_bp_debug_if = slots_4_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4768 = _T_545 ? issue_slots_4_uop_bp_debug_if : _GEN_4570; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_xcpt_ma_if = slots_4_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4769 = _T_545 ? issue_slots_4_uop_xcpt_ma_if : _GEN_4571; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_xcpt_ae_if = slots_4_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4770 = _T_545 ? issue_slots_4_uop_xcpt_ae_if : _GEN_4572; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_xcpt_pf_if = slots_4_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4771 = _T_545 ? issue_slots_4_uop_xcpt_pf_if : _GEN_4573; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_fp_single = slots_4_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4772 = _T_545 ? issue_slots_4_uop_fp_single : _GEN_4574; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_fp_val = slots_4_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4773 = _T_545 ? issue_slots_4_uop_fp_val : _GEN_4575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_frs3_en = slots_4_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4774 = _T_545 ? issue_slots_4_uop_frs3_en : _GEN_4576; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_lrs2_rtype = slots_4_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4775 = _T_545 ? issue_slots_4_uop_lrs2_rtype : _GEN_4577; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_lrs1_rtype = slots_4_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4776 = _T_545 ? issue_slots_4_uop_lrs1_rtype : _GEN_4578; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_dst_rtype = slots_4_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4777 = _T_545 ? issue_slots_4_uop_dst_rtype : _GEN_4579; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ldst_val = slots_4_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4778 = _T_545 ? issue_slots_4_uop_ldst_val : _GEN_4580; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_lrs3 = slots_4_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4779 = _T_545 ? issue_slots_4_uop_lrs3 : _GEN_4581; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_lrs2 = slots_4_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4780 = _T_545 ? issue_slots_4_uop_lrs2 : _GEN_4582; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_lrs1 = slots_4_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4781 = _T_545 ? issue_slots_4_uop_lrs1 : _GEN_4583; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_ldst = slots_4_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4782 = _T_545 ? issue_slots_4_uop_ldst : _GEN_4584; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ldst_is_rs1 = slots_4_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4783 = _T_545 ? issue_slots_4_uop_ldst_is_rs1 : _GEN_4585; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_flush_on_commit = slots_4_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4784 = _T_545 ? issue_slots_4_uop_flush_on_commit : _GEN_4586; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_unique = slots_4_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4785 = _T_545 ? issue_slots_4_uop_is_unique : _GEN_4587; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_sys_pc2epc = slots_4_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4786 = _T_545 ? issue_slots_4_uop_is_sys_pc2epc : _GEN_4588; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_uses_stq = slots_4_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4787 = _T_545 ? issue_slots_4_uop_uses_stq : _GEN_4589; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_uses_ldq = slots_4_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4788 = _T_545 ? issue_slots_4_uop_uses_ldq : _GEN_4590; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_amo = slots_4_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4789 = _T_545 ? issue_slots_4_uop_is_amo : _GEN_4591; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_fencei = slots_4_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4790 = _T_545 ? issue_slots_4_uop_is_fencei : _GEN_4592; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_fence = slots_4_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4791 = _T_545 ? issue_slots_4_uop_is_fence : _GEN_4593; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_mem_signed = slots_4_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4792 = _T_545 ? issue_slots_4_uop_mem_signed : _GEN_4594; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_mem_size = slots_4_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4793 = _T_545 ? issue_slots_4_uop_mem_size : _GEN_4595; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_mem_cmd = slots_4_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4794 = _T_545 ? issue_slots_4_uop_mem_cmd : _GEN_4596; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_bypassable = slots_4_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4795 = _T_545 ? issue_slots_4_uop_bypassable : _GEN_4597; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_4_uop_exc_cause = slots_4_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4796 = _T_545 ? issue_slots_4_uop_exc_cause : _GEN_4598; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_exception = slots_4_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4797 = _T_545 ? issue_slots_4_uop_exception : _GEN_4599; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_stale_pdst = slots_4_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4798 = _T_545 ? issue_slots_4_uop_stale_pdst : _GEN_4600; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ppred_busy = slots_4_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4799 = _T_545 ? issue_slots_4_uop_ppred_busy : _GEN_4601; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_prs3_busy = slots_4_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4800 = _T_545 ? issue_slots_4_uop_prs3_busy : _GEN_4602; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_prs2_busy = slots_4_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4801 = _T_545 ? issue_slots_4_uop_prs2_busy : _GEN_4603; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_prs1_busy = slots_4_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4802 = _T_545 ? issue_slots_4_uop_prs1_busy : _GEN_4604; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_ppred = slots_4_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4803 = _T_545 ? issue_slots_4_uop_ppred : _GEN_4605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_prs3 = slots_4_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4804 = _T_545 ? issue_slots_4_uop_prs3 : _GEN_4606; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_prs2 = slots_4_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4805 = _T_545 ? issue_slots_4_uop_prs2 : _GEN_4607; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_prs1 = slots_4_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4806 = _T_545 ? issue_slots_4_uop_prs1 : _GEN_4608; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_pdst = slots_4_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4807 = _T_545 ? issue_slots_4_uop_pdst : _GEN_4609; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_rxq_idx = slots_4_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4808 = _T_545 ? issue_slots_4_uop_rxq_idx : _GEN_4610; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_stq_idx = slots_4_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4809 = _T_545 ? issue_slots_4_uop_stq_idx : _GEN_4611; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_ldq_idx = slots_4_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4810 = _T_545 ? issue_slots_4_uop_ldq_idx : _GEN_4612; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_rob_idx = slots_4_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4811 = _T_545 ? issue_slots_4_uop_rob_idx : _GEN_4613; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_4_uop_csr_addr = slots_4_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4812 = _T_545 ? issue_slots_4_uop_csr_addr : _GEN_4614; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_4_uop_imm_packed = slots_4_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4813 = _T_545 ? issue_slots_4_uop_imm_packed : _GEN_4615; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_taken = slots_4_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4814 = _T_545 ? issue_slots_4_uop_taken : _GEN_4616; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_pc_lob = slots_4_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4815 = _T_545 ? issue_slots_4_uop_pc_lob : _GEN_4617; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_edge_inst = slots_4_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4816 = _T_545 ? issue_slots_4_uop_edge_inst : _GEN_4618; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_ftq_idx = slots_4_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4817 = _T_545 ? issue_slots_4_uop_ftq_idx : _GEN_4619; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_br_tag = slots_4_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4818 = _T_545 ? issue_slots_4_uop_br_tag : _GEN_4620; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_4_uop_br_mask = slots_4_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4819 = _T_545 ? issue_slots_4_uop_br_mask : _GEN_4621; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_sfb = slots_4_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4820 = _T_545 ? issue_slots_4_uop_is_sfb : _GEN_4622; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_jal = slots_4_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4821 = _T_545 ? issue_slots_4_uop_is_jal : _GEN_4623; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_jalr = slots_4_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4822 = _T_545 ? issue_slots_4_uop_is_jalr : _GEN_4624; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_br = slots_4_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4823 = _T_545 ? issue_slots_4_uop_is_br : _GEN_4625; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_iw_p2_poisoned = slots_4_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4824 = _T_545 ? issue_slots_4_uop_iw_p2_poisoned : _GEN_4626; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_iw_p1_poisoned = slots_4_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4825 = _T_545 ? issue_slots_4_uop_iw_p1_poisoned : _GEN_4627; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_iw_state = slots_4_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4826 = _T_545 ? issue_slots_4_uop_iw_state : _GEN_4628; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_ctrl_op3_sel = slots_4_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4827 = _T_545 ? issue_slots_4_uop_ctrl_op3_sel : _GEN_4629; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_is_std = slots_4_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4828 = _T_545 ? issue_slots_4_uop_ctrl_is_std : _GEN_4630; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_is_sta = slots_4_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4829 = _T_545 ? issue_slots_4_uop_ctrl_is_sta : _GEN_4631; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_is_load = slots_4_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4830 = _T_545 ? issue_slots_4_uop_ctrl_is_load : _GEN_4632; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_ctrl_csr_cmd = slots_4_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4831 = _T_545 ? issue_slots_4_uop_ctrl_csr_cmd : _GEN_4633; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_fcn_dw = slots_4_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4832 = _T_545 ? issue_slots_4_uop_ctrl_fcn_dw : _GEN_4634; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_ctrl_op_fcn = slots_4_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4833 = _T_545 ? issue_slots_4_uop_ctrl_op_fcn : _GEN_4635; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_ctrl_imm_sel = slots_4_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4834 = _T_545 ? issue_slots_4_uop_ctrl_imm_sel : _GEN_4636; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_ctrl_op2_sel = slots_4_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4835 = _T_545 ? issue_slots_4_uop_ctrl_op2_sel : _GEN_4637; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_ctrl_op1_sel = slots_4_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4836 = _T_545 ? issue_slots_4_uop_ctrl_op1_sel : _GEN_4638; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_ctrl_br_type = slots_4_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4837 = _T_545 ? issue_slots_4_uop_ctrl_br_type : _GEN_4639; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4838 = _T_545 ? issue_slots_4_uop_fu_code : _GEN_4640; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_iq_type = slots_4_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4839 = _T_545 ? issue_slots_4_uop_iq_type : _GEN_4641; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_4_uop_debug_pc = slots_4_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4840 = _T_545 ? issue_slots_4_uop_debug_pc : _GEN_4642; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_rvc = slots_4_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4841 = _T_545 ? issue_slots_4_uop_is_rvc : _GEN_4643; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_4_uop_debug_inst = slots_4_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4842 = _T_545 ? issue_slots_4_uop_debug_inst : _GEN_4644; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_4_uop_inst = slots_4_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4843 = _T_545 ? issue_slots_4_uop_inst : _GEN_4645; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_uopc = slots_4_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4844 = _T_545 ? issue_slots_4_uop_uopc : _GEN_4646; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_address_num = slots_4_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4845 = _T_545 ? issue_slots_4_uop_address_num : _GEN_4647; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_rob_inst_idx = slots_4_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4846 = _T_545 ? issue_slots_4_uop_rob_inst_idx : _GEN_4648; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_self_index = slots_4_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4847 = _T_545 ? issue_slots_4_uop_self_index : _GEN_4649; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_split_num = slots_4_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4848 = _T_545 ? issue_slots_4_uop_split_num : _GEN_4650; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_op2_sel = slots_4_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4849 = _T_545 ? issue_slots_4_uop_op2_sel : _GEN_4651; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_op1_sel = slots_4_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4850 = _T_545 ? issue_slots_4_uop_op1_sel : _GEN_4652; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_stale_pflag = slots_4_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4851 = _T_545 ? issue_slots_4_uop_stale_pflag : _GEN_4653; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_pflag_busy = slots_4_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4852 = _T_545 ? issue_slots_4_uop_pflag_busy : _GEN_4654; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_pwflag = slots_4_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4853 = _T_545 ? issue_slots_4_uop_pwflag : _GEN_4655; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_prflag = slots_4_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4854 = _T_545 ? issue_slots_4_uop_prflag : _GEN_4656; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_wflag = slots_4_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4855 = _T_545 ? issue_slots_4_uop_wflag : _GEN_4657; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_rflag = slots_4_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4856 = _T_545 ? issue_slots_4_uop_rflag : _GEN_4658; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_lrs3_rtype = slots_4_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4857 = _T_545 ? issue_slots_4_uop_lrs3_rtype : _GEN_4659; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_shift = slots_4_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4858 = _T_545 ? issue_slots_4_uop_shift : _GEN_4660; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_unicore = slots_4_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4859 = _T_545 ? issue_slots_4_uop_is_unicore : _GEN_4661; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_switch_off = slots_4_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4860 = _T_545 ? issue_slots_4_uop_switch_off : _GEN_4662; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_switch = slots_4_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4861 = _T_545 ? issue_slots_4_uop_switch : _GEN_4663; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4863 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 | (issue_slots_3_request & ~_T_515 & _T_518 & ~
    _T_497 | (_T_496 & ~_T_467 | (issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428)
     | issue_slots_0_request & ~_T_423 & _T_428))); // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 124:26]
  wire [1:0] _GEN_4864 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_debug_tsrc : _GEN_4666; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4865 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_debug_fsrc : _GEN_4667; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4866 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_bp_xcpt_if : _GEN_4668; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4867 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_bp_debug_if : _GEN_4669; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4868 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_xcpt_ma_if : _GEN_4670; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4869 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_xcpt_ae_if : _GEN_4671; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4870 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_xcpt_pf_if : _GEN_4672; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4871 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_fp_single : _GEN_4673; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4872 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_fp_val : _GEN_4674; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4873 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_frs3_en : _GEN_4675; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4874 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_lrs2_rtype : _GEN_4676; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4875 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_lrs1_rtype : _GEN_4677; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4876 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_dst_rtype : _GEN_4678; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4877 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ldst_val : _GEN_4679; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4878 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_lrs3 : _GEN_4680; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4879 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_lrs2 : _GEN_4681; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4880 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_lrs1 : _GEN_4682; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4881 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ldst : _GEN_4683; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4882 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ldst_is_rs1 : _GEN_4684; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4883 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_flush_on_commit : _GEN_4685; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4884 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_unique : _GEN_4686; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4885 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_sys_pc2epc : _GEN_4687; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4886 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_uses_stq : _GEN_4688; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4887 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_uses_ldq : _GEN_4689; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4888 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_amo : _GEN_4690; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4889 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_fencei : _GEN_4691; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4890 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_fence : _GEN_4692; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4891 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_mem_signed : _GEN_4693; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4892 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_mem_size : _GEN_4694; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4893 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_mem_cmd : _GEN_4695; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4894 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_bypassable : _GEN_4696; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_4895 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_exc_cause : _GEN_4697; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4896 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_exception : _GEN_4698; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4897 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_stale_pdst : _GEN_4699; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4898 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ppred_busy : _GEN_4700; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4899 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_prs3_busy : _GEN_4701; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4900 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_prs2_busy : _GEN_4702; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4901 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_prs1_busy : _GEN_4703; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4902 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ppred : _GEN_4704; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4903 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_prs3 : _GEN_4705; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4904 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_prs2 : _GEN_4706; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4905 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_prs1 : _GEN_4707; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4906 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_pdst : _GEN_4708; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4907 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_rxq_idx : _GEN_4709; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4908 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_stq_idx : _GEN_4710; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4909 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ldq_idx : _GEN_4711; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4910 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_rob_idx : _GEN_4712; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4911 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_csr_addr : _GEN_4713; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_4912 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_imm_packed : _GEN_4714; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4913 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_taken : _GEN_4715; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4914 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_pc_lob : _GEN_4716; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4915 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_edge_inst : _GEN_4717; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_4916 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ftq_idx : _GEN_4718; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4917 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_br_tag : _GEN_4719; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_4918 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_br_mask : _GEN_4720; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4919 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_sfb : _GEN_4721; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4920 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_jal : _GEN_4722; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4921 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_jalr : _GEN_4723; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4922 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_br : _GEN_4724; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4923 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_iw_p2_poisoned : _GEN_4725; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4924 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_iw_p1_poisoned : _GEN_4726; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4925 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_iw_state : _GEN_4727; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4926 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_op3_sel : _GEN_4728
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4927 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_is_std : _GEN_4729; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4928 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_is_sta : _GEN_4730; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4929 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_is_load : _GEN_4731; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4930 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_csr_cmd : _GEN_4732
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4931 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_fcn_dw : _GEN_4733; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4932 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_op_fcn : _GEN_4734; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4933 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_imm_sel : _GEN_4735
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4934 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_op2_sel : _GEN_4736
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4935 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_op1_sel : _GEN_4737
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4936 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_ctrl_br_type : _GEN_4738
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4937 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_fu_code : _GEN_4739; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4938 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_iq_type : _GEN_4740; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_4939 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_debug_pc : _GEN_4741; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4940 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_rvc : _GEN_4742; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4941 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_debug_inst : _GEN_4743; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_4942 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_inst : _GEN_4744; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_4943 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_uopc : _GEN_4745; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4944 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_address_num : _GEN_4746; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4945 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_rob_inst_idx : _GEN_4747
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4946 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_self_index : _GEN_4748; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_4947 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_split_num : _GEN_4749; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4948 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_op2_sel : _GEN_4750; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4949 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_op1_sel : _GEN_4751; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4950 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_stale_pflag : _GEN_4752; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4951 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_pflag_busy : _GEN_4753; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4952 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_pwflag : _GEN_4754; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_4953 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_prflag : _GEN_4755; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4954 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_wflag : _GEN_4756; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4955 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_rflag : _GEN_4757; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_4956 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_lrs3_rtype : _GEN_4758; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_4957 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_shift : _GEN_4759; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4958 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_is_unicore : _GEN_4760; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4959 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_switch_off : _GEN_4761; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_4960 = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 ? issue_slots_4_uop_switch : _GEN_4762; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_debug_tsrc = slots_5_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4963 = _T_575 ? issue_slots_5_uop_debug_tsrc : _GEN_4765; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_debug_fsrc = slots_5_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4964 = _T_575 ? issue_slots_5_uop_debug_fsrc : _GEN_4766; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_bp_xcpt_if = slots_5_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4965 = _T_575 ? issue_slots_5_uop_bp_xcpt_if : _GEN_4767; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_bp_debug_if = slots_5_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4966 = _T_575 ? issue_slots_5_uop_bp_debug_if : _GEN_4768; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_xcpt_ma_if = slots_5_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4967 = _T_575 ? issue_slots_5_uop_xcpt_ma_if : _GEN_4769; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_xcpt_ae_if = slots_5_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4968 = _T_575 ? issue_slots_5_uop_xcpt_ae_if : _GEN_4770; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_xcpt_pf_if = slots_5_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4969 = _T_575 ? issue_slots_5_uop_xcpt_pf_if : _GEN_4771; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_fp_single = slots_5_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4970 = _T_575 ? issue_slots_5_uop_fp_single : _GEN_4772; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_fp_val = slots_5_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4971 = _T_575 ? issue_slots_5_uop_fp_val : _GEN_4773; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_frs3_en = slots_5_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4972 = _T_575 ? issue_slots_5_uop_frs3_en : _GEN_4774; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_lrs2_rtype = slots_5_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4973 = _T_575 ? issue_slots_5_uop_lrs2_rtype : _GEN_4775; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_lrs1_rtype = slots_5_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4974 = _T_575 ? issue_slots_5_uop_lrs1_rtype : _GEN_4776; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_dst_rtype = slots_5_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4975 = _T_575 ? issue_slots_5_uop_dst_rtype : _GEN_4777; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ldst_val = slots_5_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4976 = _T_575 ? issue_slots_5_uop_ldst_val : _GEN_4778; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_lrs3 = slots_5_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4977 = _T_575 ? issue_slots_5_uop_lrs3 : _GEN_4779; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_lrs2 = slots_5_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4978 = _T_575 ? issue_slots_5_uop_lrs2 : _GEN_4780; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_lrs1 = slots_5_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4979 = _T_575 ? issue_slots_5_uop_lrs1 : _GEN_4781; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_ldst = slots_5_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4980 = _T_575 ? issue_slots_5_uop_ldst : _GEN_4782; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ldst_is_rs1 = slots_5_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4981 = _T_575 ? issue_slots_5_uop_ldst_is_rs1 : _GEN_4783; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_flush_on_commit = slots_5_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4982 = _T_575 ? issue_slots_5_uop_flush_on_commit : _GEN_4784; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_unique = slots_5_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4983 = _T_575 ? issue_slots_5_uop_is_unique : _GEN_4785; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_sys_pc2epc = slots_5_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4984 = _T_575 ? issue_slots_5_uop_is_sys_pc2epc : _GEN_4786; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_uses_stq = slots_5_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4985 = _T_575 ? issue_slots_5_uop_uses_stq : _GEN_4787; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_uses_ldq = slots_5_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4986 = _T_575 ? issue_slots_5_uop_uses_ldq : _GEN_4788; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_amo = slots_5_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4987 = _T_575 ? issue_slots_5_uop_is_amo : _GEN_4789; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_fencei = slots_5_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4988 = _T_575 ? issue_slots_5_uop_is_fencei : _GEN_4790; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_fence = slots_5_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4989 = _T_575 ? issue_slots_5_uop_is_fence : _GEN_4791; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_mem_signed = slots_5_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4990 = _T_575 ? issue_slots_5_uop_mem_signed : _GEN_4792; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_mem_size = slots_5_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4991 = _T_575 ? issue_slots_5_uop_mem_size : _GEN_4793; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_mem_cmd = slots_5_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4992 = _T_575 ? issue_slots_5_uop_mem_cmd : _GEN_4794; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_bypassable = slots_5_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4993 = _T_575 ? issue_slots_5_uop_bypassable : _GEN_4795; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_5_uop_exc_cause = slots_5_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4994 = _T_575 ? issue_slots_5_uop_exc_cause : _GEN_4796; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_exception = slots_5_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4995 = _T_575 ? issue_slots_5_uop_exception : _GEN_4797; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_stale_pdst = slots_5_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4996 = _T_575 ? issue_slots_5_uop_stale_pdst : _GEN_4798; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ppred_busy = slots_5_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4997 = _T_575 ? issue_slots_5_uop_ppred_busy : _GEN_4799; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_prs3_busy = slots_5_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4998 = _T_575 ? issue_slots_5_uop_prs3_busy : _GEN_4800; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_prs2_busy = slots_5_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4999 = _T_575 ? issue_slots_5_uop_prs2_busy : _GEN_4801; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_prs1_busy = slots_5_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5000 = _T_575 ? issue_slots_5_uop_prs1_busy : _GEN_4802; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_ppred = slots_5_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5001 = _T_575 ? issue_slots_5_uop_ppred : _GEN_4803; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_prs3 = slots_5_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5002 = _T_575 ? issue_slots_5_uop_prs3 : _GEN_4804; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_prs2 = slots_5_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5003 = _T_575 ? issue_slots_5_uop_prs2 : _GEN_4805; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_prs1 = slots_5_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5004 = _T_575 ? issue_slots_5_uop_prs1 : _GEN_4806; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_pdst = slots_5_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5005 = _T_575 ? issue_slots_5_uop_pdst : _GEN_4807; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_rxq_idx = slots_5_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5006 = _T_575 ? issue_slots_5_uop_rxq_idx : _GEN_4808; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_stq_idx = slots_5_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5007 = _T_575 ? issue_slots_5_uop_stq_idx : _GEN_4809; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_ldq_idx = slots_5_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5008 = _T_575 ? issue_slots_5_uop_ldq_idx : _GEN_4810; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_rob_idx = slots_5_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5009 = _T_575 ? issue_slots_5_uop_rob_idx : _GEN_4811; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_5_uop_csr_addr = slots_5_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5010 = _T_575 ? issue_slots_5_uop_csr_addr : _GEN_4812; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_5_uop_imm_packed = slots_5_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_5011 = _T_575 ? issue_slots_5_uop_imm_packed : _GEN_4813; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_taken = slots_5_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5012 = _T_575 ? issue_slots_5_uop_taken : _GEN_4814; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_pc_lob = slots_5_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5013 = _T_575 ? issue_slots_5_uop_pc_lob : _GEN_4815; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_edge_inst = slots_5_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5014 = _T_575 ? issue_slots_5_uop_edge_inst : _GEN_4816; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_ftq_idx = slots_5_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5015 = _T_575 ? issue_slots_5_uop_ftq_idx : _GEN_4817; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_br_tag = slots_5_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5016 = _T_575 ? issue_slots_5_uop_br_tag : _GEN_4818; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_5_uop_br_mask = slots_5_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5017 = _T_575 ? issue_slots_5_uop_br_mask : _GEN_4819; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_sfb = slots_5_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5018 = _T_575 ? issue_slots_5_uop_is_sfb : _GEN_4820; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_jal = slots_5_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5019 = _T_575 ? issue_slots_5_uop_is_jal : _GEN_4821; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_jalr = slots_5_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5020 = _T_575 ? issue_slots_5_uop_is_jalr : _GEN_4822; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_br = slots_5_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5021 = _T_575 ? issue_slots_5_uop_is_br : _GEN_4823; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_iw_p2_poisoned = slots_5_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5022 = _T_575 ? issue_slots_5_uop_iw_p2_poisoned : _GEN_4824; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_iw_p1_poisoned = slots_5_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5023 = _T_575 ? issue_slots_5_uop_iw_p1_poisoned : _GEN_4825; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_iw_state = slots_5_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5024 = _T_575 ? issue_slots_5_uop_iw_state : _GEN_4826; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_ctrl_op3_sel = slots_5_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5025 = _T_575 ? issue_slots_5_uop_ctrl_op3_sel : _GEN_4827; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_is_std = slots_5_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5026 = _T_575 ? issue_slots_5_uop_ctrl_is_std : _GEN_4828; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_is_sta = slots_5_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5027 = _T_575 ? issue_slots_5_uop_ctrl_is_sta : _GEN_4829; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_is_load = slots_5_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5028 = _T_575 ? issue_slots_5_uop_ctrl_is_load : _GEN_4830; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_ctrl_csr_cmd = slots_5_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5029 = _T_575 ? issue_slots_5_uop_ctrl_csr_cmd : _GEN_4831; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_fcn_dw = slots_5_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5030 = _T_575 ? issue_slots_5_uop_ctrl_fcn_dw : _GEN_4832; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_ctrl_op_fcn = slots_5_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5031 = _T_575 ? issue_slots_5_uop_ctrl_op_fcn : _GEN_4833; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_ctrl_imm_sel = slots_5_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5032 = _T_575 ? issue_slots_5_uop_ctrl_imm_sel : _GEN_4834; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_ctrl_op2_sel = slots_5_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5033 = _T_575 ? issue_slots_5_uop_ctrl_op2_sel : _GEN_4835; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_ctrl_op1_sel = slots_5_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5034 = _T_575 ? issue_slots_5_uop_ctrl_op1_sel : _GEN_4836; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_ctrl_br_type = slots_5_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5035 = _T_575 ? issue_slots_5_uop_ctrl_br_type : _GEN_4837; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5036 = _T_575 ? issue_slots_5_uop_fu_code : _GEN_4838; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_iq_type = slots_5_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5037 = _T_575 ? issue_slots_5_uop_iq_type : _GEN_4839; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_5_uop_debug_pc = slots_5_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_5038 = _T_575 ? issue_slots_5_uop_debug_pc : _GEN_4840; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_rvc = slots_5_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5039 = _T_575 ? issue_slots_5_uop_is_rvc : _GEN_4841; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_5_uop_debug_inst = slots_5_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5040 = _T_575 ? issue_slots_5_uop_debug_inst : _GEN_4842; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_5_uop_inst = slots_5_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5041 = _T_575 ? issue_slots_5_uop_inst : _GEN_4843; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_uopc = slots_5_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5042 = _T_575 ? issue_slots_5_uop_uopc : _GEN_4844; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_address_num = slots_5_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5043 = _T_575 ? issue_slots_5_uop_address_num : _GEN_4845; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_rob_inst_idx = slots_5_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5044 = _T_575 ? issue_slots_5_uop_rob_inst_idx : _GEN_4846; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_self_index = slots_5_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5045 = _T_575 ? issue_slots_5_uop_self_index : _GEN_4847; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_split_num = slots_5_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5046 = _T_575 ? issue_slots_5_uop_split_num : _GEN_4848; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_op2_sel = slots_5_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5047 = _T_575 ? issue_slots_5_uop_op2_sel : _GEN_4849; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_op1_sel = slots_5_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5048 = _T_575 ? issue_slots_5_uop_op1_sel : _GEN_4850; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_stale_pflag = slots_5_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5049 = _T_575 ? issue_slots_5_uop_stale_pflag : _GEN_4851; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_pflag_busy = slots_5_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5050 = _T_575 ? issue_slots_5_uop_pflag_busy : _GEN_4852; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_pwflag = slots_5_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5051 = _T_575 ? issue_slots_5_uop_pwflag : _GEN_4853; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_prflag = slots_5_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5052 = _T_575 ? issue_slots_5_uop_prflag : _GEN_4854; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_wflag = slots_5_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5053 = _T_575 ? issue_slots_5_uop_wflag : _GEN_4855; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_rflag = slots_5_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5054 = _T_575 ? issue_slots_5_uop_rflag : _GEN_4856; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_lrs3_rtype = slots_5_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5055 = _T_575 ? issue_slots_5_uop_lrs3_rtype : _GEN_4857; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_shift = slots_5_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5056 = _T_575 ? issue_slots_5_uop_shift : _GEN_4858; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_unicore = slots_5_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5057 = _T_575 ? issue_slots_5_uop_is_unicore : _GEN_4859; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_switch_off = slots_5_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5058 = _T_575 ? issue_slots_5_uop_switch_off : _GEN_4860; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_switch = slots_5_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5059 = _T_575 ? issue_slots_5_uop_switch : _GEN_4861; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5062 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_debug_tsrc : _GEN_4864; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5063 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_debug_fsrc : _GEN_4865; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5064 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_bp_xcpt_if : _GEN_4866; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5065 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_bp_debug_if : _GEN_4867; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5066 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_xcpt_ma_if : _GEN_4868; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5067 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_xcpt_ae_if : _GEN_4869; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5068 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_xcpt_pf_if : _GEN_4870; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5069 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_fp_single : _GEN_4871; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5070 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_fp_val : _GEN_4872; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5071 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_frs3_en : _GEN_4873; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5072 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_lrs2_rtype : _GEN_4874; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5073 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_lrs1_rtype : _GEN_4875; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5074 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_dst_rtype : _GEN_4876; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5075 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ldst_val : _GEN_4877; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5076 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_lrs3 : _GEN_4878; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5077 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_lrs2 : _GEN_4879; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5078 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_lrs1 : _GEN_4880; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5079 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ldst : _GEN_4881; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5080 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ldst_is_rs1 : _GEN_4882; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5081 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_flush_on_commit : _GEN_4883; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5082 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_unique : _GEN_4884; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5083 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_sys_pc2epc : _GEN_4885; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5084 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_uses_stq : _GEN_4886; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5085 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_uses_ldq : _GEN_4887; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5086 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_amo : _GEN_4888; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5087 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_fencei : _GEN_4889; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5088 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_fence : _GEN_4890; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5089 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_mem_signed : _GEN_4891; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5090 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_mem_size : _GEN_4892; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5091 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_mem_cmd : _GEN_4893; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5092 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_bypassable : _GEN_4894; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_5093 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_exc_cause : _GEN_4895; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5094 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_exception : _GEN_4896; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5095 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_stale_pdst : _GEN_4897; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5096 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ppred_busy : _GEN_4898; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5097 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_prs3_busy : _GEN_4899; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5098 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_prs2_busy : _GEN_4900; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5099 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_prs1_busy : _GEN_4901; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5100 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ppred : _GEN_4902; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5101 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_prs3 : _GEN_4903; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5102 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_prs2 : _GEN_4904; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5103 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_prs1 : _GEN_4905; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5104 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_pdst : _GEN_4906; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5105 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_rxq_idx : _GEN_4907; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5106 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_stq_idx : _GEN_4908; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5107 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ldq_idx : _GEN_4909; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5108 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_rob_idx : _GEN_4910; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5109 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_csr_addr : _GEN_4911; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_5110 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_imm_packed : _GEN_4912; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5111 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_taken : _GEN_4913; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5112 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_pc_lob : _GEN_4914; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5113 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_edge_inst : _GEN_4915; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5114 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ftq_idx : _GEN_4916; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5115 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_br_tag : _GEN_4917; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5116 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_br_mask : _GEN_4918; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5117 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_sfb : _GEN_4919; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5118 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_jal : _GEN_4920; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5119 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_jalr : _GEN_4921; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5120 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_br : _GEN_4922; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5121 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_iw_p2_poisoned : _GEN_4923; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5122 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_iw_p1_poisoned : _GEN_4924; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5123 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_iw_state : _GEN_4925; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5124 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_op3_sel : _GEN_4926
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5125 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_is_std : _GEN_4927; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5126 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_is_sta : _GEN_4928; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5127 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_is_load : _GEN_4929; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5128 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_csr_cmd : _GEN_4930
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5129 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_fcn_dw : _GEN_4931; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5130 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_op_fcn : _GEN_4932; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5131 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_imm_sel : _GEN_4933
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5132 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_op2_sel : _GEN_4934
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5133 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_op1_sel : _GEN_4935
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5134 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_ctrl_br_type : _GEN_4936
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5135 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_fu_code : _GEN_4937; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5136 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_iq_type : _GEN_4938; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_5137 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_debug_pc : _GEN_4939; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5138 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_rvc : _GEN_4940; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5139 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_debug_inst : _GEN_4941; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5140 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_inst : _GEN_4942; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5141 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_uopc : _GEN_4943; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5142 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_address_num : _GEN_4944; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5143 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_rob_inst_idx : _GEN_4945
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5144 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_self_index : _GEN_4946; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5145 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_split_num : _GEN_4947; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5146 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_op2_sel : _GEN_4948; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5147 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_op1_sel : _GEN_4949; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5148 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_stale_pflag : _GEN_4950; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5149 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_pflag_busy : _GEN_4951; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5150 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_pwflag : _GEN_4952; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5151 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_prflag : _GEN_4953; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5152 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_wflag : _GEN_4954; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5153 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_rflag : _GEN_4955; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5154 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_lrs3_rtype : _GEN_4956; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5155 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_shift : _GEN_4957; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5156 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_is_unicore : _GEN_4958; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5157 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_switch_off : _GEN_4959; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5158 = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 ? issue_slots_5_uop_switch : _GEN_4960; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_debug_tsrc = slots_6_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5161 = _T_605 ? issue_slots_6_uop_debug_tsrc : _GEN_4963; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_debug_fsrc = slots_6_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5162 = _T_605 ? issue_slots_6_uop_debug_fsrc : _GEN_4964; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_bp_xcpt_if = slots_6_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5163 = _T_605 ? issue_slots_6_uop_bp_xcpt_if : _GEN_4965; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_bp_debug_if = slots_6_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5164 = _T_605 ? issue_slots_6_uop_bp_debug_if : _GEN_4966; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_xcpt_ma_if = slots_6_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5165 = _T_605 ? issue_slots_6_uop_xcpt_ma_if : _GEN_4967; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_xcpt_ae_if = slots_6_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5166 = _T_605 ? issue_slots_6_uop_xcpt_ae_if : _GEN_4968; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_xcpt_pf_if = slots_6_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5167 = _T_605 ? issue_slots_6_uop_xcpt_pf_if : _GEN_4969; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_fp_single = slots_6_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5168 = _T_605 ? issue_slots_6_uop_fp_single : _GEN_4970; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_fp_val = slots_6_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5169 = _T_605 ? issue_slots_6_uop_fp_val : _GEN_4971; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_frs3_en = slots_6_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5170 = _T_605 ? issue_slots_6_uop_frs3_en : _GEN_4972; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_lrs2_rtype = slots_6_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5171 = _T_605 ? issue_slots_6_uop_lrs2_rtype : _GEN_4973; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_lrs1_rtype = slots_6_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5172 = _T_605 ? issue_slots_6_uop_lrs1_rtype : _GEN_4974; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_dst_rtype = slots_6_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5173 = _T_605 ? issue_slots_6_uop_dst_rtype : _GEN_4975; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ldst_val = slots_6_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5174 = _T_605 ? issue_slots_6_uop_ldst_val : _GEN_4976; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_lrs3 = slots_6_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5175 = _T_605 ? issue_slots_6_uop_lrs3 : _GEN_4977; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_lrs2 = slots_6_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5176 = _T_605 ? issue_slots_6_uop_lrs2 : _GEN_4978; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_lrs1 = slots_6_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5177 = _T_605 ? issue_slots_6_uop_lrs1 : _GEN_4979; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_ldst = slots_6_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5178 = _T_605 ? issue_slots_6_uop_ldst : _GEN_4980; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ldst_is_rs1 = slots_6_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5179 = _T_605 ? issue_slots_6_uop_ldst_is_rs1 : _GEN_4981; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_flush_on_commit = slots_6_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5180 = _T_605 ? issue_slots_6_uop_flush_on_commit : _GEN_4982; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_unique = slots_6_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5181 = _T_605 ? issue_slots_6_uop_is_unique : _GEN_4983; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_sys_pc2epc = slots_6_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5182 = _T_605 ? issue_slots_6_uop_is_sys_pc2epc : _GEN_4984; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_uses_stq = slots_6_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5183 = _T_605 ? issue_slots_6_uop_uses_stq : _GEN_4985; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_uses_ldq = slots_6_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5184 = _T_605 ? issue_slots_6_uop_uses_ldq : _GEN_4986; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_amo = slots_6_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5185 = _T_605 ? issue_slots_6_uop_is_amo : _GEN_4987; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_fencei = slots_6_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5186 = _T_605 ? issue_slots_6_uop_is_fencei : _GEN_4988; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_fence = slots_6_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5187 = _T_605 ? issue_slots_6_uop_is_fence : _GEN_4989; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_mem_signed = slots_6_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5188 = _T_605 ? issue_slots_6_uop_mem_signed : _GEN_4990; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_mem_size = slots_6_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5189 = _T_605 ? issue_slots_6_uop_mem_size : _GEN_4991; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_mem_cmd = slots_6_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5190 = _T_605 ? issue_slots_6_uop_mem_cmd : _GEN_4992; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_bypassable = slots_6_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5191 = _T_605 ? issue_slots_6_uop_bypassable : _GEN_4993; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_6_uop_exc_cause = slots_6_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_5192 = _T_605 ? issue_slots_6_uop_exc_cause : _GEN_4994; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_exception = slots_6_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5193 = _T_605 ? issue_slots_6_uop_exception : _GEN_4995; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_stale_pdst = slots_6_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5194 = _T_605 ? issue_slots_6_uop_stale_pdst : _GEN_4996; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ppred_busy = slots_6_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5195 = _T_605 ? issue_slots_6_uop_ppred_busy : _GEN_4997; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_prs3_busy = slots_6_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5196 = _T_605 ? issue_slots_6_uop_prs3_busy : _GEN_4998; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_prs2_busy = slots_6_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5197 = _T_605 ? issue_slots_6_uop_prs2_busy : _GEN_4999; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_prs1_busy = slots_6_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5198 = _T_605 ? issue_slots_6_uop_prs1_busy : _GEN_5000; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_ppred = slots_6_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5199 = _T_605 ? issue_slots_6_uop_ppred : _GEN_5001; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_prs3 = slots_6_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5200 = _T_605 ? issue_slots_6_uop_prs3 : _GEN_5002; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_prs2 = slots_6_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5201 = _T_605 ? issue_slots_6_uop_prs2 : _GEN_5003; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_prs1 = slots_6_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5202 = _T_605 ? issue_slots_6_uop_prs1 : _GEN_5004; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_pdst = slots_6_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5203 = _T_605 ? issue_slots_6_uop_pdst : _GEN_5005; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_rxq_idx = slots_6_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5204 = _T_605 ? issue_slots_6_uop_rxq_idx : _GEN_5006; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_stq_idx = slots_6_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5205 = _T_605 ? issue_slots_6_uop_stq_idx : _GEN_5007; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_ldq_idx = slots_6_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5206 = _T_605 ? issue_slots_6_uop_ldq_idx : _GEN_5008; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_rob_idx = slots_6_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5207 = _T_605 ? issue_slots_6_uop_rob_idx : _GEN_5009; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_6_uop_csr_addr = slots_6_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5208 = _T_605 ? issue_slots_6_uop_csr_addr : _GEN_5010; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_6_uop_imm_packed = slots_6_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_5209 = _T_605 ? issue_slots_6_uop_imm_packed : _GEN_5011; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_taken = slots_6_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5210 = _T_605 ? issue_slots_6_uop_taken : _GEN_5012; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_pc_lob = slots_6_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5211 = _T_605 ? issue_slots_6_uop_pc_lob : _GEN_5013; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_edge_inst = slots_6_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5212 = _T_605 ? issue_slots_6_uop_edge_inst : _GEN_5014; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_ftq_idx = slots_6_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5213 = _T_605 ? issue_slots_6_uop_ftq_idx : _GEN_5015; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_br_tag = slots_6_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5214 = _T_605 ? issue_slots_6_uop_br_tag : _GEN_5016; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_6_uop_br_mask = slots_6_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5215 = _T_605 ? issue_slots_6_uop_br_mask : _GEN_5017; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_sfb = slots_6_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5216 = _T_605 ? issue_slots_6_uop_is_sfb : _GEN_5018; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_jal = slots_6_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5217 = _T_605 ? issue_slots_6_uop_is_jal : _GEN_5019; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_jalr = slots_6_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5218 = _T_605 ? issue_slots_6_uop_is_jalr : _GEN_5020; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_br = slots_6_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5219 = _T_605 ? issue_slots_6_uop_is_br : _GEN_5021; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_iw_p2_poisoned = slots_6_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5220 = _T_605 ? issue_slots_6_uop_iw_p2_poisoned : _GEN_5022; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_iw_p1_poisoned = slots_6_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5221 = _T_605 ? issue_slots_6_uop_iw_p1_poisoned : _GEN_5023; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_iw_state = slots_6_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5222 = _T_605 ? issue_slots_6_uop_iw_state : _GEN_5024; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_ctrl_op3_sel = slots_6_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5223 = _T_605 ? issue_slots_6_uop_ctrl_op3_sel : _GEN_5025; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_is_std = slots_6_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5224 = _T_605 ? issue_slots_6_uop_ctrl_is_std : _GEN_5026; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_is_sta = slots_6_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5225 = _T_605 ? issue_slots_6_uop_ctrl_is_sta : _GEN_5027; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_is_load = slots_6_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5226 = _T_605 ? issue_slots_6_uop_ctrl_is_load : _GEN_5028; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_ctrl_csr_cmd = slots_6_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5227 = _T_605 ? issue_slots_6_uop_ctrl_csr_cmd : _GEN_5029; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_fcn_dw = slots_6_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5228 = _T_605 ? issue_slots_6_uop_ctrl_fcn_dw : _GEN_5030; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_ctrl_op_fcn = slots_6_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5229 = _T_605 ? issue_slots_6_uop_ctrl_op_fcn : _GEN_5031; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_ctrl_imm_sel = slots_6_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5230 = _T_605 ? issue_slots_6_uop_ctrl_imm_sel : _GEN_5032; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_ctrl_op2_sel = slots_6_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5231 = _T_605 ? issue_slots_6_uop_ctrl_op2_sel : _GEN_5033; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_ctrl_op1_sel = slots_6_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5232 = _T_605 ? issue_slots_6_uop_ctrl_op1_sel : _GEN_5034; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_ctrl_br_type = slots_6_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5233 = _T_605 ? issue_slots_6_uop_ctrl_br_type : _GEN_5035; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5234 = _T_605 ? issue_slots_6_uop_fu_code : _GEN_5036; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_iq_type = slots_6_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5235 = _T_605 ? issue_slots_6_uop_iq_type : _GEN_5037; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_6_uop_debug_pc = slots_6_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_5236 = _T_605 ? issue_slots_6_uop_debug_pc : _GEN_5038; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_rvc = slots_6_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5237 = _T_605 ? issue_slots_6_uop_is_rvc : _GEN_5039; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_6_uop_debug_inst = slots_6_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5238 = _T_605 ? issue_slots_6_uop_debug_inst : _GEN_5040; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_6_uop_inst = slots_6_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5239 = _T_605 ? issue_slots_6_uop_inst : _GEN_5041; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_uopc = slots_6_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5240 = _T_605 ? issue_slots_6_uop_uopc : _GEN_5042; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_address_num = slots_6_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5241 = _T_605 ? issue_slots_6_uop_address_num : _GEN_5043; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_rob_inst_idx = slots_6_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5242 = _T_605 ? issue_slots_6_uop_rob_inst_idx : _GEN_5044; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_self_index = slots_6_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5243 = _T_605 ? issue_slots_6_uop_self_index : _GEN_5045; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_split_num = slots_6_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5244 = _T_605 ? issue_slots_6_uop_split_num : _GEN_5046; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_op2_sel = slots_6_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5245 = _T_605 ? issue_slots_6_uop_op2_sel : _GEN_5047; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_op1_sel = slots_6_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5246 = _T_605 ? issue_slots_6_uop_op1_sel : _GEN_5048; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_stale_pflag = slots_6_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5247 = _T_605 ? issue_slots_6_uop_stale_pflag : _GEN_5049; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_pflag_busy = slots_6_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5248 = _T_605 ? issue_slots_6_uop_pflag_busy : _GEN_5050; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_pwflag = slots_6_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5249 = _T_605 ? issue_slots_6_uop_pwflag : _GEN_5051; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_prflag = slots_6_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5250 = _T_605 ? issue_slots_6_uop_prflag : _GEN_5052; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_wflag = slots_6_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5251 = _T_605 ? issue_slots_6_uop_wflag : _GEN_5053; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_rflag = slots_6_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5252 = _T_605 ? issue_slots_6_uop_rflag : _GEN_5054; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_lrs3_rtype = slots_6_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5253 = _T_605 ? issue_slots_6_uop_lrs3_rtype : _GEN_5055; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_shift = slots_6_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5254 = _T_605 ? issue_slots_6_uop_shift : _GEN_5056; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_unicore = slots_6_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5255 = _T_605 ? issue_slots_6_uop_is_unicore : _GEN_5057; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_switch_off = slots_6_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5256 = _T_605 ? issue_slots_6_uop_switch_off : _GEN_5058; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_switch = slots_6_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5257 = _T_605 ? issue_slots_6_uop_switch : _GEN_5059; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5260 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_debug_tsrc : _GEN_5062; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5261 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_debug_fsrc : _GEN_5063; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5262 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_bp_xcpt_if : _GEN_5064; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5263 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_bp_debug_if : _GEN_5065; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5264 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_xcpt_ma_if : _GEN_5066; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5265 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_xcpt_ae_if : _GEN_5067; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5266 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_xcpt_pf_if : _GEN_5068; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5267 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_fp_single : _GEN_5069; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5268 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_fp_val : _GEN_5070; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5269 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_frs3_en : _GEN_5071; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5270 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_lrs2_rtype : _GEN_5072; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5271 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_lrs1_rtype : _GEN_5073; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5272 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_dst_rtype : _GEN_5074; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5273 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ldst_val : _GEN_5075; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5274 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_lrs3 : _GEN_5076; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5275 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_lrs2 : _GEN_5077; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5276 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_lrs1 : _GEN_5078; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5277 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ldst : _GEN_5079; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5278 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ldst_is_rs1 : _GEN_5080; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5279 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_flush_on_commit : _GEN_5081; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5280 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_unique : _GEN_5082; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5281 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_sys_pc2epc : _GEN_5083; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5282 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_uses_stq : _GEN_5084; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5283 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_uses_ldq : _GEN_5085; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5284 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_amo : _GEN_5086; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5285 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_fencei : _GEN_5087; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5286 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_fence : _GEN_5088; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5287 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_mem_signed : _GEN_5089; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5288 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_mem_size : _GEN_5090; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5289 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_mem_cmd : _GEN_5091; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5290 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_bypassable : _GEN_5092; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_5291 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_exc_cause : _GEN_5093; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5292 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_exception : _GEN_5094; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5293 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_stale_pdst : _GEN_5095; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5294 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ppred_busy : _GEN_5096; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5295 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_prs3_busy : _GEN_5097; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5296 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_prs2_busy : _GEN_5098; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5297 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_prs1_busy : _GEN_5099; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5298 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ppred : _GEN_5100; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5299 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_prs3 : _GEN_5101; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5300 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_prs2 : _GEN_5102; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5301 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_prs1 : _GEN_5103; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5302 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_pdst : _GEN_5104; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5303 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_rxq_idx : _GEN_5105; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5304 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_stq_idx : _GEN_5106; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5305 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ldq_idx : _GEN_5107; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5306 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_rob_idx : _GEN_5108; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5307 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_csr_addr : _GEN_5109; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_5308 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_imm_packed : _GEN_5110; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5309 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_taken : _GEN_5111; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5310 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_pc_lob : _GEN_5112; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5311 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_edge_inst : _GEN_5113; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5312 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ftq_idx : _GEN_5114; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5313 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_br_tag : _GEN_5115; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5314 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_br_mask : _GEN_5116; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5315 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_sfb : _GEN_5117; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5316 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_jal : _GEN_5118; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5317 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_jalr : _GEN_5119; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5318 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_br : _GEN_5120; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5319 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_iw_p2_poisoned : _GEN_5121; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5320 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_iw_p1_poisoned : _GEN_5122; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5321 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_iw_state : _GEN_5123; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5322 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_op3_sel : _GEN_5124
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5323 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_is_std : _GEN_5125; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5324 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_is_sta : _GEN_5126; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5325 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_is_load : _GEN_5127; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5326 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_csr_cmd : _GEN_5128
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5327 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_fcn_dw : _GEN_5129; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5328 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_op_fcn : _GEN_5130; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5329 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_imm_sel : _GEN_5131
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5330 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_op2_sel : _GEN_5132
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5331 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_op1_sel : _GEN_5133
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5332 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_ctrl_br_type : _GEN_5134
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5333 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_fu_code : _GEN_5135; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5334 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_iq_type : _GEN_5136; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_5335 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_debug_pc : _GEN_5137; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5336 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_rvc : _GEN_5138; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5337 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_debug_inst : _GEN_5139; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5338 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_inst : _GEN_5140; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5339 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_uopc : _GEN_5141; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5340 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_address_num : _GEN_5142; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5341 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_rob_inst_idx : _GEN_5143
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5342 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_self_index : _GEN_5144; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5343 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_split_num : _GEN_5145; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5344 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_op2_sel : _GEN_5146; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5345 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_op1_sel : _GEN_5147; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5346 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_stale_pflag : _GEN_5148; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5347 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_pflag_busy : _GEN_5149; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5348 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_pwflag : _GEN_5150; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5349 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_prflag : _GEN_5151; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5350 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_wflag : _GEN_5152; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5351 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_rflag : _GEN_5153; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5352 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_lrs3_rtype : _GEN_5154; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5353 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_shift : _GEN_5155; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5354 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_is_unicore : _GEN_5156; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5355 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_switch_off : _GEN_5157; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5356 = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 ? issue_slots_6_uop_switch : _GEN_5158; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_debug_tsrc = slots_7_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5359 = _T_635 ? issue_slots_7_uop_debug_tsrc : _GEN_5161; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_debug_fsrc = slots_7_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5360 = _T_635 ? issue_slots_7_uop_debug_fsrc : _GEN_5162; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_bp_xcpt_if = slots_7_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5361 = _T_635 ? issue_slots_7_uop_bp_xcpt_if : _GEN_5163; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_bp_debug_if = slots_7_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5362 = _T_635 ? issue_slots_7_uop_bp_debug_if : _GEN_5164; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_xcpt_ma_if = slots_7_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5363 = _T_635 ? issue_slots_7_uop_xcpt_ma_if : _GEN_5165; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_xcpt_ae_if = slots_7_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5364 = _T_635 ? issue_slots_7_uop_xcpt_ae_if : _GEN_5166; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_xcpt_pf_if = slots_7_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5365 = _T_635 ? issue_slots_7_uop_xcpt_pf_if : _GEN_5167; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_fp_single = slots_7_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5366 = _T_635 ? issue_slots_7_uop_fp_single : _GEN_5168; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_fp_val = slots_7_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5367 = _T_635 ? issue_slots_7_uop_fp_val : _GEN_5169; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_frs3_en = slots_7_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5368 = _T_635 ? issue_slots_7_uop_frs3_en : _GEN_5170; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_lrs2_rtype = slots_7_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5369 = _T_635 ? issue_slots_7_uop_lrs2_rtype : _GEN_5171; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_lrs1_rtype = slots_7_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5370 = _T_635 ? issue_slots_7_uop_lrs1_rtype : _GEN_5172; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_dst_rtype = slots_7_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5371 = _T_635 ? issue_slots_7_uop_dst_rtype : _GEN_5173; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ldst_val = slots_7_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5372 = _T_635 ? issue_slots_7_uop_ldst_val : _GEN_5174; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_lrs3 = slots_7_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5373 = _T_635 ? issue_slots_7_uop_lrs3 : _GEN_5175; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_lrs2 = slots_7_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5374 = _T_635 ? issue_slots_7_uop_lrs2 : _GEN_5176; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_lrs1 = slots_7_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5375 = _T_635 ? issue_slots_7_uop_lrs1 : _GEN_5177; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_ldst = slots_7_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5376 = _T_635 ? issue_slots_7_uop_ldst : _GEN_5178; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ldst_is_rs1 = slots_7_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5377 = _T_635 ? issue_slots_7_uop_ldst_is_rs1 : _GEN_5179; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_flush_on_commit = slots_7_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5378 = _T_635 ? issue_slots_7_uop_flush_on_commit : _GEN_5180; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_unique = slots_7_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5379 = _T_635 ? issue_slots_7_uop_is_unique : _GEN_5181; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_sys_pc2epc = slots_7_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5380 = _T_635 ? issue_slots_7_uop_is_sys_pc2epc : _GEN_5182; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_uses_stq = slots_7_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5381 = _T_635 ? issue_slots_7_uop_uses_stq : _GEN_5183; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_uses_ldq = slots_7_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5382 = _T_635 ? issue_slots_7_uop_uses_ldq : _GEN_5184; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_amo = slots_7_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5383 = _T_635 ? issue_slots_7_uop_is_amo : _GEN_5185; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_fencei = slots_7_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5384 = _T_635 ? issue_slots_7_uop_is_fencei : _GEN_5186; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_fence = slots_7_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5385 = _T_635 ? issue_slots_7_uop_is_fence : _GEN_5187; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_mem_signed = slots_7_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5386 = _T_635 ? issue_slots_7_uop_mem_signed : _GEN_5188; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_mem_size = slots_7_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5387 = _T_635 ? issue_slots_7_uop_mem_size : _GEN_5189; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_mem_cmd = slots_7_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5388 = _T_635 ? issue_slots_7_uop_mem_cmd : _GEN_5190; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_bypassable = slots_7_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5389 = _T_635 ? issue_slots_7_uop_bypassable : _GEN_5191; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_7_uop_exc_cause = slots_7_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_5390 = _T_635 ? issue_slots_7_uop_exc_cause : _GEN_5192; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_exception = slots_7_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5391 = _T_635 ? issue_slots_7_uop_exception : _GEN_5193; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_stale_pdst = slots_7_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5392 = _T_635 ? issue_slots_7_uop_stale_pdst : _GEN_5194; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ppred_busy = slots_7_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5393 = _T_635 ? issue_slots_7_uop_ppred_busy : _GEN_5195; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_prs3_busy = slots_7_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5394 = _T_635 ? issue_slots_7_uop_prs3_busy : _GEN_5196; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_prs2_busy = slots_7_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5395 = _T_635 ? issue_slots_7_uop_prs2_busy : _GEN_5197; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_prs1_busy = slots_7_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5396 = _T_635 ? issue_slots_7_uop_prs1_busy : _GEN_5198; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_ppred = slots_7_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5397 = _T_635 ? issue_slots_7_uop_ppred : _GEN_5199; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_prs3 = slots_7_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5398 = _T_635 ? issue_slots_7_uop_prs3 : _GEN_5200; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_prs2 = slots_7_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5399 = _T_635 ? issue_slots_7_uop_prs2 : _GEN_5201; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_prs1 = slots_7_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5400 = _T_635 ? issue_slots_7_uop_prs1 : _GEN_5202; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_pdst = slots_7_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5401 = _T_635 ? issue_slots_7_uop_pdst : _GEN_5203; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_rxq_idx = slots_7_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5402 = _T_635 ? issue_slots_7_uop_rxq_idx : _GEN_5204; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_stq_idx = slots_7_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5403 = _T_635 ? issue_slots_7_uop_stq_idx : _GEN_5205; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_ldq_idx = slots_7_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5404 = _T_635 ? issue_slots_7_uop_ldq_idx : _GEN_5206; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_rob_idx = slots_7_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5405 = _T_635 ? issue_slots_7_uop_rob_idx : _GEN_5207; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_7_uop_csr_addr = slots_7_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5406 = _T_635 ? issue_slots_7_uop_csr_addr : _GEN_5208; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_7_uop_imm_packed = slots_7_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_5407 = _T_635 ? issue_slots_7_uop_imm_packed : _GEN_5209; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_taken = slots_7_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5408 = _T_635 ? issue_slots_7_uop_taken : _GEN_5210; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_pc_lob = slots_7_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5409 = _T_635 ? issue_slots_7_uop_pc_lob : _GEN_5211; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_edge_inst = slots_7_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5410 = _T_635 ? issue_slots_7_uop_edge_inst : _GEN_5212; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_ftq_idx = slots_7_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5411 = _T_635 ? issue_slots_7_uop_ftq_idx : _GEN_5213; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_br_tag = slots_7_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5412 = _T_635 ? issue_slots_7_uop_br_tag : _GEN_5214; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_7_uop_br_mask = slots_7_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5413 = _T_635 ? issue_slots_7_uop_br_mask : _GEN_5215; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_sfb = slots_7_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5414 = _T_635 ? issue_slots_7_uop_is_sfb : _GEN_5216; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_jal = slots_7_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5415 = _T_635 ? issue_slots_7_uop_is_jal : _GEN_5217; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_jalr = slots_7_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5416 = _T_635 ? issue_slots_7_uop_is_jalr : _GEN_5218; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_br = slots_7_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5417 = _T_635 ? issue_slots_7_uop_is_br : _GEN_5219; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_iw_p2_poisoned = slots_7_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5418 = _T_635 ? issue_slots_7_uop_iw_p2_poisoned : _GEN_5220; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_iw_p1_poisoned = slots_7_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5419 = _T_635 ? issue_slots_7_uop_iw_p1_poisoned : _GEN_5221; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_iw_state = slots_7_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5420 = _T_635 ? issue_slots_7_uop_iw_state : _GEN_5222; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_ctrl_op3_sel = slots_7_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5421 = _T_635 ? issue_slots_7_uop_ctrl_op3_sel : _GEN_5223; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_is_std = slots_7_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5422 = _T_635 ? issue_slots_7_uop_ctrl_is_std : _GEN_5224; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_is_sta = slots_7_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5423 = _T_635 ? issue_slots_7_uop_ctrl_is_sta : _GEN_5225; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_is_load = slots_7_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5424 = _T_635 ? issue_slots_7_uop_ctrl_is_load : _GEN_5226; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_ctrl_csr_cmd = slots_7_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5425 = _T_635 ? issue_slots_7_uop_ctrl_csr_cmd : _GEN_5227; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_fcn_dw = slots_7_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5426 = _T_635 ? issue_slots_7_uop_ctrl_fcn_dw : _GEN_5228; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_ctrl_op_fcn = slots_7_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5427 = _T_635 ? issue_slots_7_uop_ctrl_op_fcn : _GEN_5229; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_ctrl_imm_sel = slots_7_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5428 = _T_635 ? issue_slots_7_uop_ctrl_imm_sel : _GEN_5230; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_ctrl_op2_sel = slots_7_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5429 = _T_635 ? issue_slots_7_uop_ctrl_op2_sel : _GEN_5231; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_ctrl_op1_sel = slots_7_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5430 = _T_635 ? issue_slots_7_uop_ctrl_op1_sel : _GEN_5232; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_ctrl_br_type = slots_7_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5431 = _T_635 ? issue_slots_7_uop_ctrl_br_type : _GEN_5233; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5432 = _T_635 ? issue_slots_7_uop_fu_code : _GEN_5234; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_iq_type = slots_7_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5433 = _T_635 ? issue_slots_7_uop_iq_type : _GEN_5235; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_7_uop_debug_pc = slots_7_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_5434 = _T_635 ? issue_slots_7_uop_debug_pc : _GEN_5236; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_rvc = slots_7_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5435 = _T_635 ? issue_slots_7_uop_is_rvc : _GEN_5237; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_7_uop_debug_inst = slots_7_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5436 = _T_635 ? issue_slots_7_uop_debug_inst : _GEN_5238; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_7_uop_inst = slots_7_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5437 = _T_635 ? issue_slots_7_uop_inst : _GEN_5239; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_uopc = slots_7_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5438 = _T_635 ? issue_slots_7_uop_uopc : _GEN_5240; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_address_num = slots_7_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5439 = _T_635 ? issue_slots_7_uop_address_num : _GEN_5241; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_rob_inst_idx = slots_7_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5440 = _T_635 ? issue_slots_7_uop_rob_inst_idx : _GEN_5242; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_self_index = slots_7_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5441 = _T_635 ? issue_slots_7_uop_self_index : _GEN_5243; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_split_num = slots_7_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5442 = _T_635 ? issue_slots_7_uop_split_num : _GEN_5244; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_op2_sel = slots_7_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5443 = _T_635 ? issue_slots_7_uop_op2_sel : _GEN_5245; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_op1_sel = slots_7_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5444 = _T_635 ? issue_slots_7_uop_op1_sel : _GEN_5246; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_stale_pflag = slots_7_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5445 = _T_635 ? issue_slots_7_uop_stale_pflag : _GEN_5247; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_pflag_busy = slots_7_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5446 = _T_635 ? issue_slots_7_uop_pflag_busy : _GEN_5248; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_pwflag = slots_7_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5447 = _T_635 ? issue_slots_7_uop_pwflag : _GEN_5249; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_prflag = slots_7_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5448 = _T_635 ? issue_slots_7_uop_prflag : _GEN_5250; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_wflag = slots_7_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5449 = _T_635 ? issue_slots_7_uop_wflag : _GEN_5251; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_rflag = slots_7_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5450 = _T_635 ? issue_slots_7_uop_rflag : _GEN_5252; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_lrs3_rtype = slots_7_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5451 = _T_635 ? issue_slots_7_uop_lrs3_rtype : _GEN_5253; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_shift = slots_7_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5452 = _T_635 ? issue_slots_7_uop_shift : _GEN_5254; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_unicore = slots_7_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5453 = _T_635 ? issue_slots_7_uop_is_unicore : _GEN_5255; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_switch_off = slots_7_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5454 = _T_635 ? issue_slots_7_uop_switch_off : _GEN_5256; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_switch = slots_7_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5455 = _T_635 ? issue_slots_7_uop_switch : _GEN_5257; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5458 = _T_646 & ~_T_617 ? issue_slots_7_uop_debug_tsrc : _GEN_5260; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5459 = _T_646 & ~_T_617 ? issue_slots_7_uop_debug_fsrc : _GEN_5261; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5460 = _T_646 & ~_T_617 ? issue_slots_7_uop_bp_xcpt_if : _GEN_5262; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5461 = _T_646 & ~_T_617 ? issue_slots_7_uop_bp_debug_if : _GEN_5263; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5462 = _T_646 & ~_T_617 ? issue_slots_7_uop_xcpt_ma_if : _GEN_5264; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5463 = _T_646 & ~_T_617 ? issue_slots_7_uop_xcpt_ae_if : _GEN_5265; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5464 = _T_646 & ~_T_617 ? issue_slots_7_uop_xcpt_pf_if : _GEN_5266; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5465 = _T_646 & ~_T_617 ? issue_slots_7_uop_fp_single : _GEN_5267; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5466 = _T_646 & ~_T_617 ? issue_slots_7_uop_fp_val : _GEN_5268; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5467 = _T_646 & ~_T_617 ? issue_slots_7_uop_frs3_en : _GEN_5269; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5468 = _T_646 & ~_T_617 ? issue_slots_7_uop_lrs2_rtype : _GEN_5270; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5469 = _T_646 & ~_T_617 ? issue_slots_7_uop_lrs1_rtype : _GEN_5271; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5470 = _T_646 & ~_T_617 ? issue_slots_7_uop_dst_rtype : _GEN_5272; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5471 = _T_646 & ~_T_617 ? issue_slots_7_uop_ldst_val : _GEN_5273; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5472 = _T_646 & ~_T_617 ? issue_slots_7_uop_lrs3 : _GEN_5274; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5473 = _T_646 & ~_T_617 ? issue_slots_7_uop_lrs2 : _GEN_5275; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5474 = _T_646 & ~_T_617 ? issue_slots_7_uop_lrs1 : _GEN_5276; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5475 = _T_646 & ~_T_617 ? issue_slots_7_uop_ldst : _GEN_5277; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5476 = _T_646 & ~_T_617 ? issue_slots_7_uop_ldst_is_rs1 : _GEN_5278; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5477 = _T_646 & ~_T_617 ? issue_slots_7_uop_flush_on_commit : _GEN_5279; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5478 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_unique : _GEN_5280; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5479 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_sys_pc2epc : _GEN_5281; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5480 = _T_646 & ~_T_617 ? issue_slots_7_uop_uses_stq : _GEN_5282; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5481 = _T_646 & ~_T_617 ? issue_slots_7_uop_uses_ldq : _GEN_5283; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5482 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_amo : _GEN_5284; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5483 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_fencei : _GEN_5285; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5484 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_fence : _GEN_5286; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5485 = _T_646 & ~_T_617 ? issue_slots_7_uop_mem_signed : _GEN_5287; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5486 = _T_646 & ~_T_617 ? issue_slots_7_uop_mem_size : _GEN_5288; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5487 = _T_646 & ~_T_617 ? issue_slots_7_uop_mem_cmd : _GEN_5289; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5488 = _T_646 & ~_T_617 ? issue_slots_7_uop_bypassable : _GEN_5290; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_5489 = _T_646 & ~_T_617 ? issue_slots_7_uop_exc_cause : _GEN_5291; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5490 = _T_646 & ~_T_617 ? issue_slots_7_uop_exception : _GEN_5292; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5491 = _T_646 & ~_T_617 ? issue_slots_7_uop_stale_pdst : _GEN_5293; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5492 = _T_646 & ~_T_617 ? issue_slots_7_uop_ppred_busy : _GEN_5294; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5493 = _T_646 & ~_T_617 ? issue_slots_7_uop_prs3_busy : _GEN_5295; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5494 = _T_646 & ~_T_617 ? issue_slots_7_uop_prs2_busy : _GEN_5296; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5495 = _T_646 & ~_T_617 ? issue_slots_7_uop_prs1_busy : _GEN_5297; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5496 = _T_646 & ~_T_617 ? issue_slots_7_uop_ppred : _GEN_5298; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5497 = _T_646 & ~_T_617 ? issue_slots_7_uop_prs3 : _GEN_5299; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5498 = _T_646 & ~_T_617 ? issue_slots_7_uop_prs2 : _GEN_5300; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5499 = _T_646 & ~_T_617 ? issue_slots_7_uop_prs1 : _GEN_5301; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5500 = _T_646 & ~_T_617 ? issue_slots_7_uop_pdst : _GEN_5302; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5501 = _T_646 & ~_T_617 ? issue_slots_7_uop_rxq_idx : _GEN_5303; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5502 = _T_646 & ~_T_617 ? issue_slots_7_uop_stq_idx : _GEN_5304; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5503 = _T_646 & ~_T_617 ? issue_slots_7_uop_ldq_idx : _GEN_5305; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5504 = _T_646 & ~_T_617 ? issue_slots_7_uop_rob_idx : _GEN_5306; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5505 = _T_646 & ~_T_617 ? issue_slots_7_uop_csr_addr : _GEN_5307; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_5506 = _T_646 & ~_T_617 ? issue_slots_7_uop_imm_packed : _GEN_5308; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5507 = _T_646 & ~_T_617 ? issue_slots_7_uop_taken : _GEN_5309; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5508 = _T_646 & ~_T_617 ? issue_slots_7_uop_pc_lob : _GEN_5310; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5509 = _T_646 & ~_T_617 ? issue_slots_7_uop_edge_inst : _GEN_5311; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5510 = _T_646 & ~_T_617 ? issue_slots_7_uop_ftq_idx : _GEN_5312; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5511 = _T_646 & ~_T_617 ? issue_slots_7_uop_br_tag : _GEN_5313; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5512 = _T_646 & ~_T_617 ? issue_slots_7_uop_br_mask : _GEN_5314; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5513 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_sfb : _GEN_5315; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5514 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_jal : _GEN_5316; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5515 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_jalr : _GEN_5317; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5516 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_br : _GEN_5318; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5517 = _T_646 & ~_T_617 ? issue_slots_7_uop_iw_p2_poisoned : _GEN_5319; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5518 = _T_646 & ~_T_617 ? issue_slots_7_uop_iw_p1_poisoned : _GEN_5320; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5519 = _T_646 & ~_T_617 ? issue_slots_7_uop_iw_state : _GEN_5321; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5520 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_op3_sel : _GEN_5322; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5521 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_is_std : _GEN_5323; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5522 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_is_sta : _GEN_5324; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5523 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_is_load : _GEN_5325; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5524 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_csr_cmd : _GEN_5326; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5525 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_fcn_dw : _GEN_5327; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5526 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_op_fcn : _GEN_5328; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5527 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_imm_sel : _GEN_5329; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5528 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_op2_sel : _GEN_5330; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5529 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_op1_sel : _GEN_5331; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5530 = _T_646 & ~_T_617 ? issue_slots_7_uop_ctrl_br_type : _GEN_5332; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5531 = _T_646 & ~_T_617 ? issue_slots_7_uop_fu_code : _GEN_5333; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5532 = _T_646 & ~_T_617 ? issue_slots_7_uop_iq_type : _GEN_5334; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_5533 = _T_646 & ~_T_617 ? issue_slots_7_uop_debug_pc : _GEN_5335; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5534 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_rvc : _GEN_5336; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5535 = _T_646 & ~_T_617 ? issue_slots_7_uop_debug_inst : _GEN_5337; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5536 = _T_646 & ~_T_617 ? issue_slots_7_uop_inst : _GEN_5338; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5537 = _T_646 & ~_T_617 ? issue_slots_7_uop_uopc : _GEN_5339; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5538 = _T_646 & ~_T_617 ? issue_slots_7_uop_address_num : _GEN_5340; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5539 = _T_646 & ~_T_617 ? issue_slots_7_uop_rob_inst_idx : _GEN_5341; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5540 = _T_646 & ~_T_617 ? issue_slots_7_uop_self_index : _GEN_5342; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5541 = _T_646 & ~_T_617 ? issue_slots_7_uop_split_num : _GEN_5343; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5542 = _T_646 & ~_T_617 ? issue_slots_7_uop_op2_sel : _GEN_5344; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5543 = _T_646 & ~_T_617 ? issue_slots_7_uop_op1_sel : _GEN_5345; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5544 = _T_646 & ~_T_617 ? issue_slots_7_uop_stale_pflag : _GEN_5346; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5545 = _T_646 & ~_T_617 ? issue_slots_7_uop_pflag_busy : _GEN_5347; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5546 = _T_646 & ~_T_617 ? issue_slots_7_uop_pwflag : _GEN_5348; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5547 = _T_646 & ~_T_617 ? issue_slots_7_uop_prflag : _GEN_5349; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5548 = _T_646 & ~_T_617 ? issue_slots_7_uop_wflag : _GEN_5350; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5549 = _T_646 & ~_T_617 ? issue_slots_7_uop_rflag : _GEN_5351; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5550 = _T_646 & ~_T_617 ? issue_slots_7_uop_lrs3_rtype : _GEN_5352; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5551 = _T_646 & ~_T_617 ? issue_slots_7_uop_shift : _GEN_5353; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5552 = _T_646 & ~_T_617 ? issue_slots_7_uop_is_unicore : _GEN_5354; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5553 = _T_646 & ~_T_617 ? issue_slots_7_uop_switch_off : _GEN_5355; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5554 = _T_646 & ~_T_617 ? issue_slots_7_uop_switch : _GEN_5356; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_debug_tsrc = slots_8_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5557 = _T_665 ? issue_slots_8_uop_debug_tsrc : _GEN_5359; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_debug_fsrc = slots_8_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5558 = _T_665 ? issue_slots_8_uop_debug_fsrc : _GEN_5360; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_bp_xcpt_if = slots_8_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5559 = _T_665 ? issue_slots_8_uop_bp_xcpt_if : _GEN_5361; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_bp_debug_if = slots_8_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5560 = _T_665 ? issue_slots_8_uop_bp_debug_if : _GEN_5362; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_xcpt_ma_if = slots_8_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5561 = _T_665 ? issue_slots_8_uop_xcpt_ma_if : _GEN_5363; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_xcpt_ae_if = slots_8_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5562 = _T_665 ? issue_slots_8_uop_xcpt_ae_if : _GEN_5364; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_xcpt_pf_if = slots_8_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5563 = _T_665 ? issue_slots_8_uop_xcpt_pf_if : _GEN_5365; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_fp_single = slots_8_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5564 = _T_665 ? issue_slots_8_uop_fp_single : _GEN_5366; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_fp_val = slots_8_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5565 = _T_665 ? issue_slots_8_uop_fp_val : _GEN_5367; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_frs3_en = slots_8_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5566 = _T_665 ? issue_slots_8_uop_frs3_en : _GEN_5368; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_lrs2_rtype = slots_8_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5567 = _T_665 ? issue_slots_8_uop_lrs2_rtype : _GEN_5369; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_lrs1_rtype = slots_8_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5568 = _T_665 ? issue_slots_8_uop_lrs1_rtype : _GEN_5370; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_dst_rtype = slots_8_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5569 = _T_665 ? issue_slots_8_uop_dst_rtype : _GEN_5371; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ldst_val = slots_8_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5570 = _T_665 ? issue_slots_8_uop_ldst_val : _GEN_5372; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_lrs3 = slots_8_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5571 = _T_665 ? issue_slots_8_uop_lrs3 : _GEN_5373; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_lrs2 = slots_8_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5572 = _T_665 ? issue_slots_8_uop_lrs2 : _GEN_5374; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_lrs1 = slots_8_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5573 = _T_665 ? issue_slots_8_uop_lrs1 : _GEN_5375; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_ldst = slots_8_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5574 = _T_665 ? issue_slots_8_uop_ldst : _GEN_5376; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ldst_is_rs1 = slots_8_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5575 = _T_665 ? issue_slots_8_uop_ldst_is_rs1 : _GEN_5377; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_flush_on_commit = slots_8_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5576 = _T_665 ? issue_slots_8_uop_flush_on_commit : _GEN_5378; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_unique = slots_8_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5577 = _T_665 ? issue_slots_8_uop_is_unique : _GEN_5379; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_sys_pc2epc = slots_8_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5578 = _T_665 ? issue_slots_8_uop_is_sys_pc2epc : _GEN_5380; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_uses_stq = slots_8_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5579 = _T_665 ? issue_slots_8_uop_uses_stq : _GEN_5381; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_uses_ldq = slots_8_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5580 = _T_665 ? issue_slots_8_uop_uses_ldq : _GEN_5382; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_amo = slots_8_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5581 = _T_665 ? issue_slots_8_uop_is_amo : _GEN_5383; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_fencei = slots_8_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5582 = _T_665 ? issue_slots_8_uop_is_fencei : _GEN_5384; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_fence = slots_8_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5583 = _T_665 ? issue_slots_8_uop_is_fence : _GEN_5385; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_mem_signed = slots_8_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5584 = _T_665 ? issue_slots_8_uop_mem_signed : _GEN_5386; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_mem_size = slots_8_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5585 = _T_665 ? issue_slots_8_uop_mem_size : _GEN_5387; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_mem_cmd = slots_8_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5586 = _T_665 ? issue_slots_8_uop_mem_cmd : _GEN_5388; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_bypassable = slots_8_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5587 = _T_665 ? issue_slots_8_uop_bypassable : _GEN_5389; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_8_uop_exc_cause = slots_8_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_5588 = _T_665 ? issue_slots_8_uop_exc_cause : _GEN_5390; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_exception = slots_8_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5589 = _T_665 ? issue_slots_8_uop_exception : _GEN_5391; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_stale_pdst = slots_8_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5590 = _T_665 ? issue_slots_8_uop_stale_pdst : _GEN_5392; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ppred_busy = slots_8_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5591 = _T_665 ? issue_slots_8_uop_ppred_busy : _GEN_5393; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_prs3_busy = slots_8_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5592 = _T_665 ? issue_slots_8_uop_prs3_busy : _GEN_5394; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_prs2_busy = slots_8_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5593 = _T_665 ? issue_slots_8_uop_prs2_busy : _GEN_5395; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_prs1_busy = slots_8_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5594 = _T_665 ? issue_slots_8_uop_prs1_busy : _GEN_5396; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_ppred = slots_8_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5595 = _T_665 ? issue_slots_8_uop_ppred : _GEN_5397; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_prs3 = slots_8_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5596 = _T_665 ? issue_slots_8_uop_prs3 : _GEN_5398; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_prs2 = slots_8_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5597 = _T_665 ? issue_slots_8_uop_prs2 : _GEN_5399; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_prs1 = slots_8_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5598 = _T_665 ? issue_slots_8_uop_prs1 : _GEN_5400; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_pdst = slots_8_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5599 = _T_665 ? issue_slots_8_uop_pdst : _GEN_5401; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_rxq_idx = slots_8_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5600 = _T_665 ? issue_slots_8_uop_rxq_idx : _GEN_5402; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_stq_idx = slots_8_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5601 = _T_665 ? issue_slots_8_uop_stq_idx : _GEN_5403; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_ldq_idx = slots_8_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5602 = _T_665 ? issue_slots_8_uop_ldq_idx : _GEN_5404; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_rob_idx = slots_8_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5603 = _T_665 ? issue_slots_8_uop_rob_idx : _GEN_5405; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_8_uop_csr_addr = slots_8_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5604 = _T_665 ? issue_slots_8_uop_csr_addr : _GEN_5406; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_8_uop_imm_packed = slots_8_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_5605 = _T_665 ? issue_slots_8_uop_imm_packed : _GEN_5407; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_taken = slots_8_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5606 = _T_665 ? issue_slots_8_uop_taken : _GEN_5408; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_pc_lob = slots_8_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5607 = _T_665 ? issue_slots_8_uop_pc_lob : _GEN_5409; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_edge_inst = slots_8_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5608 = _T_665 ? issue_slots_8_uop_edge_inst : _GEN_5410; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_ftq_idx = slots_8_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5609 = _T_665 ? issue_slots_8_uop_ftq_idx : _GEN_5411; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_br_tag = slots_8_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5610 = _T_665 ? issue_slots_8_uop_br_tag : _GEN_5412; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_8_uop_br_mask = slots_8_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5611 = _T_665 ? issue_slots_8_uop_br_mask : _GEN_5413; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_sfb = slots_8_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5612 = _T_665 ? issue_slots_8_uop_is_sfb : _GEN_5414; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_jal = slots_8_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5613 = _T_665 ? issue_slots_8_uop_is_jal : _GEN_5415; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_jalr = slots_8_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5614 = _T_665 ? issue_slots_8_uop_is_jalr : _GEN_5416; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_br = slots_8_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5615 = _T_665 ? issue_slots_8_uop_is_br : _GEN_5417; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_iw_p2_poisoned = slots_8_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5616 = _T_665 ? issue_slots_8_uop_iw_p2_poisoned : _GEN_5418; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_iw_p1_poisoned = slots_8_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5617 = _T_665 ? issue_slots_8_uop_iw_p1_poisoned : _GEN_5419; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_iw_state = slots_8_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5618 = _T_665 ? issue_slots_8_uop_iw_state : _GEN_5420; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_ctrl_op3_sel = slots_8_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5619 = _T_665 ? issue_slots_8_uop_ctrl_op3_sel : _GEN_5421; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_is_std = slots_8_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5620 = _T_665 ? issue_slots_8_uop_ctrl_is_std : _GEN_5422; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_is_sta = slots_8_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5621 = _T_665 ? issue_slots_8_uop_ctrl_is_sta : _GEN_5423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_is_load = slots_8_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5622 = _T_665 ? issue_slots_8_uop_ctrl_is_load : _GEN_5424; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_ctrl_csr_cmd = slots_8_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5623 = _T_665 ? issue_slots_8_uop_ctrl_csr_cmd : _GEN_5425; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_fcn_dw = slots_8_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5624 = _T_665 ? issue_slots_8_uop_ctrl_fcn_dw : _GEN_5426; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_ctrl_op_fcn = slots_8_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5625 = _T_665 ? issue_slots_8_uop_ctrl_op_fcn : _GEN_5427; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_ctrl_imm_sel = slots_8_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5626 = _T_665 ? issue_slots_8_uop_ctrl_imm_sel : _GEN_5428; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_ctrl_op2_sel = slots_8_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5627 = _T_665 ? issue_slots_8_uop_ctrl_op2_sel : _GEN_5429; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_ctrl_op1_sel = slots_8_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5628 = _T_665 ? issue_slots_8_uop_ctrl_op1_sel : _GEN_5430; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_ctrl_br_type = slots_8_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5629 = _T_665 ? issue_slots_8_uop_ctrl_br_type : _GEN_5431; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5630 = _T_665 ? issue_slots_8_uop_fu_code : _GEN_5432; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_iq_type = slots_8_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5631 = _T_665 ? issue_slots_8_uop_iq_type : _GEN_5433; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_8_uop_debug_pc = slots_8_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_5632 = _T_665 ? issue_slots_8_uop_debug_pc : _GEN_5434; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_rvc = slots_8_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5633 = _T_665 ? issue_slots_8_uop_is_rvc : _GEN_5435; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_8_uop_debug_inst = slots_8_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5634 = _T_665 ? issue_slots_8_uop_debug_inst : _GEN_5436; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_8_uop_inst = slots_8_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5635 = _T_665 ? issue_slots_8_uop_inst : _GEN_5437; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_uopc = slots_8_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5636 = _T_665 ? issue_slots_8_uop_uopc : _GEN_5438; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_address_num = slots_8_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5637 = _T_665 ? issue_slots_8_uop_address_num : _GEN_5439; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_rob_inst_idx = slots_8_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5638 = _T_665 ? issue_slots_8_uop_rob_inst_idx : _GEN_5440; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_self_index = slots_8_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5639 = _T_665 ? issue_slots_8_uop_self_index : _GEN_5441; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_split_num = slots_8_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5640 = _T_665 ? issue_slots_8_uop_split_num : _GEN_5442; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_op2_sel = slots_8_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5641 = _T_665 ? issue_slots_8_uop_op2_sel : _GEN_5443; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_op1_sel = slots_8_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5642 = _T_665 ? issue_slots_8_uop_op1_sel : _GEN_5444; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_stale_pflag = slots_8_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5643 = _T_665 ? issue_slots_8_uop_stale_pflag : _GEN_5445; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_pflag_busy = slots_8_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5644 = _T_665 ? issue_slots_8_uop_pflag_busy : _GEN_5446; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_pwflag = slots_8_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5645 = _T_665 ? issue_slots_8_uop_pwflag : _GEN_5447; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_prflag = slots_8_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5646 = _T_665 ? issue_slots_8_uop_prflag : _GEN_5448; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_wflag = slots_8_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5647 = _T_665 ? issue_slots_8_uop_wflag : _GEN_5449; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_rflag = slots_8_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5648 = _T_665 ? issue_slots_8_uop_rflag : _GEN_5450; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_lrs3_rtype = slots_8_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5649 = _T_665 ? issue_slots_8_uop_lrs3_rtype : _GEN_5451; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_shift = slots_8_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5650 = _T_665 ? issue_slots_8_uop_shift : _GEN_5452; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_unicore = slots_8_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5651 = _T_665 ? issue_slots_8_uop_is_unicore : _GEN_5453; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_switch_off = slots_8_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5652 = _T_665 ? issue_slots_8_uop_switch_off : _GEN_5454; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_switch = slots_8_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5653 = _T_665 ? issue_slots_8_uop_switch : _GEN_5455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5656 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_debug_tsrc : _GEN_5458; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5657 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_debug_fsrc : _GEN_5459; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5658 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_bp_xcpt_if : _GEN_5460; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5659 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_bp_debug_if : _GEN_5461; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5660 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_xcpt_ma_if : _GEN_5462; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5661 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_xcpt_ae_if : _GEN_5463; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5662 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_xcpt_pf_if : _GEN_5464; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5663 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_fp_single : _GEN_5465; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5664 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_fp_val : _GEN_5466; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5665 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_frs3_en : _GEN_5467; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5666 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_lrs2_rtype : _GEN_5468; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5667 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_lrs1_rtype : _GEN_5469; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5668 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_dst_rtype : _GEN_5470; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5669 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ldst_val : _GEN_5471; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5670 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_lrs3 : _GEN_5472; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5671 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_lrs2 : _GEN_5473; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5672 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_lrs1 : _GEN_5474; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5673 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ldst : _GEN_5475; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5674 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ldst_is_rs1 : _GEN_5476; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5675 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_flush_on_commit : _GEN_5477; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5676 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_unique : _GEN_5478; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5677 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_sys_pc2epc : _GEN_5479; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5678 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_uses_stq : _GEN_5480; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5679 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_uses_ldq : _GEN_5481; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5680 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_amo : _GEN_5482; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5681 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_fencei : _GEN_5483; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5682 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_fence : _GEN_5484; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5683 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_mem_signed : _GEN_5485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5684 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_mem_size : _GEN_5486; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5685 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_mem_cmd : _GEN_5487; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5686 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_bypassable : _GEN_5488; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_5687 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_exc_cause : _GEN_5489; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5688 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_exception : _GEN_5490; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5689 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_stale_pdst : _GEN_5491; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5690 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ppred_busy : _GEN_5492; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5691 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_prs3_busy : _GEN_5493; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5692 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_prs2_busy : _GEN_5494; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5693 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_prs1_busy : _GEN_5495; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5694 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ppred : _GEN_5496; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5695 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_prs3 : _GEN_5497; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5696 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_prs2 : _GEN_5498; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5697 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_prs1 : _GEN_5499; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5698 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_pdst : _GEN_5500; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5699 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_rxq_idx : _GEN_5501; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5700 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_stq_idx : _GEN_5502; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5701 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ldq_idx : _GEN_5503; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5702 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_rob_idx : _GEN_5504; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5703 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_csr_addr : _GEN_5505; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_5704 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_imm_packed : _GEN_5506; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5705 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_taken : _GEN_5507; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5706 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_pc_lob : _GEN_5508; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5707 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_edge_inst : _GEN_5509; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5708 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ftq_idx : _GEN_5510; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5709 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_br_tag : _GEN_5511; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5710 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_br_mask : _GEN_5512; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5711 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_sfb : _GEN_5513; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5712 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_jal : _GEN_5514; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5713 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_jalr : _GEN_5515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5714 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_br : _GEN_5516; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5715 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_iw_p2_poisoned : _GEN_5517; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5716 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_iw_p1_poisoned : _GEN_5518; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5717 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_iw_state : _GEN_5519; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5718 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_op3_sel : _GEN_5520
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5719 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_is_std : _GEN_5521; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5720 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_is_sta : _GEN_5522; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5721 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_is_load : _GEN_5523; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5722 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_csr_cmd : _GEN_5524
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5723 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_fcn_dw : _GEN_5525; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5724 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_op_fcn : _GEN_5526; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5725 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_imm_sel : _GEN_5527
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5726 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_op2_sel : _GEN_5528
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5727 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_op1_sel : _GEN_5529
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5728 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_ctrl_br_type : _GEN_5530
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5729 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_fu_code : _GEN_5531; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5730 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_iq_type : _GEN_5532; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_5731 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_debug_pc : _GEN_5533; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5732 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_rvc : _GEN_5534; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5733 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_debug_inst : _GEN_5535; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5734 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_inst : _GEN_5536; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5735 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_uopc : _GEN_5537; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5736 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_address_num : _GEN_5538; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5737 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_rob_inst_idx : _GEN_5539
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5738 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_self_index : _GEN_5540; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5739 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_split_num : _GEN_5541; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5740 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_op2_sel : _GEN_5542; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5741 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_op1_sel : _GEN_5543; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5742 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_stale_pflag : _GEN_5544; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5743 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_pflag_busy : _GEN_5545; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5744 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_pwflag : _GEN_5546; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5745 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_prflag : _GEN_5547; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5746 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_wflag : _GEN_5548; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5747 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_rflag : _GEN_5549; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5748 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_lrs3_rtype : _GEN_5550; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5749 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_shift : _GEN_5551; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5750 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_is_unicore : _GEN_5552; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5751 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_switch_off : _GEN_5553; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5752 = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 ? issue_slots_8_uop_switch : _GEN_5554; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_debug_tsrc = slots_9_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5755 = _T_695 ? issue_slots_9_uop_debug_tsrc : _GEN_5557; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_debug_fsrc = slots_9_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5756 = _T_695 ? issue_slots_9_uop_debug_fsrc : _GEN_5558; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_bp_xcpt_if = slots_9_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5757 = _T_695 ? issue_slots_9_uop_bp_xcpt_if : _GEN_5559; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_bp_debug_if = slots_9_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5758 = _T_695 ? issue_slots_9_uop_bp_debug_if : _GEN_5560; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_xcpt_ma_if = slots_9_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5759 = _T_695 ? issue_slots_9_uop_xcpt_ma_if : _GEN_5561; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_xcpt_ae_if = slots_9_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5760 = _T_695 ? issue_slots_9_uop_xcpt_ae_if : _GEN_5562; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_xcpt_pf_if = slots_9_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5761 = _T_695 ? issue_slots_9_uop_xcpt_pf_if : _GEN_5563; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_fp_single = slots_9_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5762 = _T_695 ? issue_slots_9_uop_fp_single : _GEN_5564; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_fp_val = slots_9_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5763 = _T_695 ? issue_slots_9_uop_fp_val : _GEN_5565; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_frs3_en = slots_9_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5764 = _T_695 ? issue_slots_9_uop_frs3_en : _GEN_5566; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_lrs2_rtype = slots_9_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5765 = _T_695 ? issue_slots_9_uop_lrs2_rtype : _GEN_5567; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_lrs1_rtype = slots_9_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5766 = _T_695 ? issue_slots_9_uop_lrs1_rtype : _GEN_5568; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_dst_rtype = slots_9_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5767 = _T_695 ? issue_slots_9_uop_dst_rtype : _GEN_5569; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ldst_val = slots_9_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5768 = _T_695 ? issue_slots_9_uop_ldst_val : _GEN_5570; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_lrs3 = slots_9_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5769 = _T_695 ? issue_slots_9_uop_lrs3 : _GEN_5571; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_lrs2 = slots_9_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5770 = _T_695 ? issue_slots_9_uop_lrs2 : _GEN_5572; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_lrs1 = slots_9_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5771 = _T_695 ? issue_slots_9_uop_lrs1 : _GEN_5573; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_ldst = slots_9_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5772 = _T_695 ? issue_slots_9_uop_ldst : _GEN_5574; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ldst_is_rs1 = slots_9_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5773 = _T_695 ? issue_slots_9_uop_ldst_is_rs1 : _GEN_5575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_flush_on_commit = slots_9_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5774 = _T_695 ? issue_slots_9_uop_flush_on_commit : _GEN_5576; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_unique = slots_9_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5775 = _T_695 ? issue_slots_9_uop_is_unique : _GEN_5577; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_sys_pc2epc = slots_9_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5776 = _T_695 ? issue_slots_9_uop_is_sys_pc2epc : _GEN_5578; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_uses_stq = slots_9_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5777 = _T_695 ? issue_slots_9_uop_uses_stq : _GEN_5579; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_uses_ldq = slots_9_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5778 = _T_695 ? issue_slots_9_uop_uses_ldq : _GEN_5580; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_amo = slots_9_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5779 = _T_695 ? issue_slots_9_uop_is_amo : _GEN_5581; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_fencei = slots_9_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5780 = _T_695 ? issue_slots_9_uop_is_fencei : _GEN_5582; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_fence = slots_9_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5781 = _T_695 ? issue_slots_9_uop_is_fence : _GEN_5583; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_mem_signed = slots_9_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5782 = _T_695 ? issue_slots_9_uop_mem_signed : _GEN_5584; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_mem_size = slots_9_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5783 = _T_695 ? issue_slots_9_uop_mem_size : _GEN_5585; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_mem_cmd = slots_9_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5784 = _T_695 ? issue_slots_9_uop_mem_cmd : _GEN_5586; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_bypassable = slots_9_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5785 = _T_695 ? issue_slots_9_uop_bypassable : _GEN_5587; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_9_uop_exc_cause = slots_9_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_5786 = _T_695 ? issue_slots_9_uop_exc_cause : _GEN_5588; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_exception = slots_9_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5787 = _T_695 ? issue_slots_9_uop_exception : _GEN_5589; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_stale_pdst = slots_9_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5788 = _T_695 ? issue_slots_9_uop_stale_pdst : _GEN_5590; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ppred_busy = slots_9_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5789 = _T_695 ? issue_slots_9_uop_ppred_busy : _GEN_5591; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_prs3_busy = slots_9_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5790 = _T_695 ? issue_slots_9_uop_prs3_busy : _GEN_5592; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_prs2_busy = slots_9_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5791 = _T_695 ? issue_slots_9_uop_prs2_busy : _GEN_5593; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_prs1_busy = slots_9_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5792 = _T_695 ? issue_slots_9_uop_prs1_busy : _GEN_5594; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_ppred = slots_9_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5793 = _T_695 ? issue_slots_9_uop_ppred : _GEN_5595; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_prs3 = slots_9_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5794 = _T_695 ? issue_slots_9_uop_prs3 : _GEN_5596; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_prs2 = slots_9_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5795 = _T_695 ? issue_slots_9_uop_prs2 : _GEN_5597; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_prs1 = slots_9_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5796 = _T_695 ? issue_slots_9_uop_prs1 : _GEN_5598; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_pdst = slots_9_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5797 = _T_695 ? issue_slots_9_uop_pdst : _GEN_5599; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_rxq_idx = slots_9_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5798 = _T_695 ? issue_slots_9_uop_rxq_idx : _GEN_5600; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_stq_idx = slots_9_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5799 = _T_695 ? issue_slots_9_uop_stq_idx : _GEN_5601; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_ldq_idx = slots_9_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5800 = _T_695 ? issue_slots_9_uop_ldq_idx : _GEN_5602; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_rob_idx = slots_9_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5801 = _T_695 ? issue_slots_9_uop_rob_idx : _GEN_5603; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_9_uop_csr_addr = slots_9_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5802 = _T_695 ? issue_slots_9_uop_csr_addr : _GEN_5604; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_9_uop_imm_packed = slots_9_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_5803 = _T_695 ? issue_slots_9_uop_imm_packed : _GEN_5605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_taken = slots_9_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5804 = _T_695 ? issue_slots_9_uop_taken : _GEN_5606; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_pc_lob = slots_9_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5805 = _T_695 ? issue_slots_9_uop_pc_lob : _GEN_5607; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_edge_inst = slots_9_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5806 = _T_695 ? issue_slots_9_uop_edge_inst : _GEN_5608; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_ftq_idx = slots_9_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5807 = _T_695 ? issue_slots_9_uop_ftq_idx : _GEN_5609; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_br_tag = slots_9_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5808 = _T_695 ? issue_slots_9_uop_br_tag : _GEN_5610; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_9_uop_br_mask = slots_9_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_5809 = _T_695 ? issue_slots_9_uop_br_mask : _GEN_5611; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_sfb = slots_9_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5810 = _T_695 ? issue_slots_9_uop_is_sfb : _GEN_5612; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_jal = slots_9_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5811 = _T_695 ? issue_slots_9_uop_is_jal : _GEN_5613; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_jalr = slots_9_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5812 = _T_695 ? issue_slots_9_uop_is_jalr : _GEN_5614; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_br = slots_9_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5813 = _T_695 ? issue_slots_9_uop_is_br : _GEN_5615; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_iw_p2_poisoned = slots_9_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5814 = _T_695 ? issue_slots_9_uop_iw_p2_poisoned : _GEN_5616; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_iw_p1_poisoned = slots_9_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5815 = _T_695 ? issue_slots_9_uop_iw_p1_poisoned : _GEN_5617; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_iw_state = slots_9_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5816 = _T_695 ? issue_slots_9_uop_iw_state : _GEN_5618; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_ctrl_op3_sel = slots_9_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5817 = _T_695 ? issue_slots_9_uop_ctrl_op3_sel : _GEN_5619; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_is_std = slots_9_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5818 = _T_695 ? issue_slots_9_uop_ctrl_is_std : _GEN_5620; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_is_sta = slots_9_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5819 = _T_695 ? issue_slots_9_uop_ctrl_is_sta : _GEN_5621; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_is_load = slots_9_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5820 = _T_695 ? issue_slots_9_uop_ctrl_is_load : _GEN_5622; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_ctrl_csr_cmd = slots_9_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5821 = _T_695 ? issue_slots_9_uop_ctrl_csr_cmd : _GEN_5623; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_fcn_dw = slots_9_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5822 = _T_695 ? issue_slots_9_uop_ctrl_fcn_dw : _GEN_5624; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_ctrl_op_fcn = slots_9_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5823 = _T_695 ? issue_slots_9_uop_ctrl_op_fcn : _GEN_5625; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_ctrl_imm_sel = slots_9_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5824 = _T_695 ? issue_slots_9_uop_ctrl_imm_sel : _GEN_5626; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_ctrl_op2_sel = slots_9_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5825 = _T_695 ? issue_slots_9_uop_ctrl_op2_sel : _GEN_5627; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_ctrl_op1_sel = slots_9_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5826 = _T_695 ? issue_slots_9_uop_ctrl_op1_sel : _GEN_5628; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_ctrl_br_type = slots_9_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5827 = _T_695 ? issue_slots_9_uop_ctrl_br_type : _GEN_5629; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5828 = _T_695 ? issue_slots_9_uop_fu_code : _GEN_5630; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_iq_type = slots_9_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5829 = _T_695 ? issue_slots_9_uop_iq_type : _GEN_5631; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_9_uop_debug_pc = slots_9_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_5830 = _T_695 ? issue_slots_9_uop_debug_pc : _GEN_5632; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_rvc = slots_9_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5831 = _T_695 ? issue_slots_9_uop_is_rvc : _GEN_5633; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_9_uop_debug_inst = slots_9_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5832 = _T_695 ? issue_slots_9_uop_debug_inst : _GEN_5634; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_9_uop_inst = slots_9_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_5833 = _T_695 ? issue_slots_9_uop_inst : _GEN_5635; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_uopc = slots_9_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5834 = _T_695 ? issue_slots_9_uop_uopc : _GEN_5636; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_address_num = slots_9_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5835 = _T_695 ? issue_slots_9_uop_address_num : _GEN_5637; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_rob_inst_idx = slots_9_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5836 = _T_695 ? issue_slots_9_uop_rob_inst_idx : _GEN_5638; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_self_index = slots_9_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5837 = _T_695 ? issue_slots_9_uop_self_index : _GEN_5639; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_split_num = slots_9_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5838 = _T_695 ? issue_slots_9_uop_split_num : _GEN_5640; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_op2_sel = slots_9_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5839 = _T_695 ? issue_slots_9_uop_op2_sel : _GEN_5641; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_op1_sel = slots_9_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5840 = _T_695 ? issue_slots_9_uop_op1_sel : _GEN_5642; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_stale_pflag = slots_9_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5841 = _T_695 ? issue_slots_9_uop_stale_pflag : _GEN_5643; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_pflag_busy = slots_9_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5842 = _T_695 ? issue_slots_9_uop_pflag_busy : _GEN_5644; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_pwflag = slots_9_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5843 = _T_695 ? issue_slots_9_uop_pwflag : _GEN_5645; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_prflag = slots_9_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_5844 = _T_695 ? issue_slots_9_uop_prflag : _GEN_5646; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_wflag = slots_9_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5845 = _T_695 ? issue_slots_9_uop_wflag : _GEN_5647; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_rflag = slots_9_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5846 = _T_695 ? issue_slots_9_uop_rflag : _GEN_5648; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_lrs3_rtype = slots_9_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5847 = _T_695 ? issue_slots_9_uop_lrs3_rtype : _GEN_5649; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_shift = slots_9_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_5848 = _T_695 ? issue_slots_9_uop_shift : _GEN_5650; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_unicore = slots_9_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5849 = _T_695 ? issue_slots_9_uop_is_unicore : _GEN_5651; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_switch_off = slots_9_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5850 = _T_695 ? issue_slots_9_uop_switch_off : _GEN_5652; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_switch = slots_9_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5851 = _T_695 ? issue_slots_9_uop_switch : _GEN_5653; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5853 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 | (issue_slots_8_request & ~_T_665 & _T_668 & ~
    _T_647 | (_T_646 & ~_T_617 | (issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 | (issue_slots_5_request & ~_T_575
     & _T_578 & ~_T_557 | _GEN_4863)))); // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 124:26]
  wire [1:0] _GEN_5854 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_debug_tsrc : _GEN_5656; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5855 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_debug_fsrc : _GEN_5657; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5856 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_bp_xcpt_if : _GEN_5658; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5857 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_bp_debug_if : _GEN_5659; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5858 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_xcpt_ma_if : _GEN_5660; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5859 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_xcpt_ae_if : _GEN_5661; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5860 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_xcpt_pf_if : _GEN_5662; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5861 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_fp_single : _GEN_5663; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5862 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_fp_val : _GEN_5664; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5863 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_frs3_en : _GEN_5665; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5864 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_lrs2_rtype : _GEN_5666; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5865 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_lrs1_rtype : _GEN_5667; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5866 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_dst_rtype : _GEN_5668; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5867 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ldst_val : _GEN_5669; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5868 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_lrs3 : _GEN_5670; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5869 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_lrs2 : _GEN_5671; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5870 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_lrs1 : _GEN_5672; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5871 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ldst : _GEN_5673; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5872 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ldst_is_rs1 : _GEN_5674; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5873 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_flush_on_commit : _GEN_5675; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5874 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_unique : _GEN_5676; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5875 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_sys_pc2epc : _GEN_5677; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5876 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_uses_stq : _GEN_5678; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5877 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_uses_ldq : _GEN_5679; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5878 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_amo : _GEN_5680; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5879 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_fencei : _GEN_5681; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5880 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_fence : _GEN_5682; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5881 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_mem_signed : _GEN_5683; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5882 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_mem_size : _GEN_5684; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5883 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_mem_cmd : _GEN_5685; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5884 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_bypassable : _GEN_5686; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_5885 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_exc_cause : _GEN_5687; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5886 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_exception : _GEN_5688; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5887 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_stale_pdst : _GEN_5689; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5888 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ppred_busy : _GEN_5690; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5889 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_prs3_busy : _GEN_5691; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5890 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_prs2_busy : _GEN_5692; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5891 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_prs1_busy : _GEN_5693; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5892 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ppred : _GEN_5694; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5893 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_prs3 : _GEN_5695; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5894 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_prs2 : _GEN_5696; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5895 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_prs1 : _GEN_5697; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5896 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_pdst : _GEN_5698; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5897 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_rxq_idx : _GEN_5699; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5898 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_stq_idx : _GEN_5700; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5899 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ldq_idx : _GEN_5701; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5900 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_rob_idx : _GEN_5702; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5901 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_csr_addr : _GEN_5703; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_5902 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_imm_packed : _GEN_5704; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5903 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_taken : _GEN_5705; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5904 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_pc_lob : _GEN_5706; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5905 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_edge_inst : _GEN_5707; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_5906 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ftq_idx : _GEN_5708; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5907 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_br_tag : _GEN_5709; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_5908 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_br_mask : _GEN_5710; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5909 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_sfb : _GEN_5711; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5910 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_jal : _GEN_5712; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5911 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_jalr : _GEN_5713; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5912 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_br : _GEN_5714; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5913 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_iw_p2_poisoned : _GEN_5715; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5914 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_iw_p1_poisoned : _GEN_5716; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5915 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_iw_state : _GEN_5717; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5916 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_op3_sel : _GEN_5718
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5917 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_is_std : _GEN_5719; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5918 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_is_sta : _GEN_5720; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5919 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_is_load : _GEN_5721; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5920 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_csr_cmd : _GEN_5722
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5921 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_fcn_dw : _GEN_5723; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5922 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_op_fcn : _GEN_5724; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5923 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_imm_sel : _GEN_5725
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5924 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_op2_sel : _GEN_5726
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5925 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_op1_sel : _GEN_5727
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5926 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_ctrl_br_type : _GEN_5728
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_5927 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_fu_code : _GEN_5729; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5928 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_iq_type : _GEN_5730; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_5929 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_debug_pc : _GEN_5731; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5930 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_rvc : _GEN_5732; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5931 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_debug_inst : _GEN_5733; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_5932 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_inst : _GEN_5734; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_5933 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_uopc : _GEN_5735; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5934 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_address_num : _GEN_5736; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5935 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_rob_inst_idx : _GEN_5737
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5936 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_self_index : _GEN_5738; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_5937 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_split_num : _GEN_5739; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5938 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_op2_sel : _GEN_5740; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5939 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_op1_sel : _GEN_5741; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5940 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_stale_pflag : _GEN_5742; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5941 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_pflag_busy : _GEN_5743; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5942 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_pwflag : _GEN_5744; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_5943 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_prflag : _GEN_5745; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5944 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_wflag : _GEN_5746; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5945 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_rflag : _GEN_5747; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_5946 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_lrs3_rtype : _GEN_5748; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_5947 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_shift : _GEN_5749; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5948 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_is_unicore : _GEN_5750; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5949 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_switch_off : _GEN_5751; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_5950 = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 ? issue_slots_9_uop_switch : _GEN_5752; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_debug_tsrc = slots_10_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5953 = _T_725 ? issue_slots_10_uop_debug_tsrc : _GEN_5755; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_debug_fsrc = slots_10_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5954 = _T_725 ? issue_slots_10_uop_debug_fsrc : _GEN_5756; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_bp_xcpt_if = slots_10_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5955 = _T_725 ? issue_slots_10_uop_bp_xcpt_if : _GEN_5757; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_bp_debug_if = slots_10_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5956 = _T_725 ? issue_slots_10_uop_bp_debug_if : _GEN_5758; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_xcpt_ma_if = slots_10_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5957 = _T_725 ? issue_slots_10_uop_xcpt_ma_if : _GEN_5759; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_xcpt_ae_if = slots_10_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5958 = _T_725 ? issue_slots_10_uop_xcpt_ae_if : _GEN_5760; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_xcpt_pf_if = slots_10_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5959 = _T_725 ? issue_slots_10_uop_xcpt_pf_if : _GEN_5761; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_fp_single = slots_10_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5960 = _T_725 ? issue_slots_10_uop_fp_single : _GEN_5762; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_fp_val = slots_10_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5961 = _T_725 ? issue_slots_10_uop_fp_val : _GEN_5763; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_frs3_en = slots_10_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5962 = _T_725 ? issue_slots_10_uop_frs3_en : _GEN_5764; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_lrs2_rtype = slots_10_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5963 = _T_725 ? issue_slots_10_uop_lrs2_rtype : _GEN_5765; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_lrs1_rtype = slots_10_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5964 = _T_725 ? issue_slots_10_uop_lrs1_rtype : _GEN_5766; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_dst_rtype = slots_10_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5965 = _T_725 ? issue_slots_10_uop_dst_rtype : _GEN_5767; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ldst_val = slots_10_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5966 = _T_725 ? issue_slots_10_uop_ldst_val : _GEN_5768; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_lrs3 = slots_10_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5967 = _T_725 ? issue_slots_10_uop_lrs3 : _GEN_5769; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_lrs2 = slots_10_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5968 = _T_725 ? issue_slots_10_uop_lrs2 : _GEN_5770; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_lrs1 = slots_10_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5969 = _T_725 ? issue_slots_10_uop_lrs1 : _GEN_5771; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_ldst = slots_10_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5970 = _T_725 ? issue_slots_10_uop_ldst : _GEN_5772; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ldst_is_rs1 = slots_10_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5971 = _T_725 ? issue_slots_10_uop_ldst_is_rs1 : _GEN_5773; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_flush_on_commit = slots_10_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5972 = _T_725 ? issue_slots_10_uop_flush_on_commit : _GEN_5774; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_unique = slots_10_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5973 = _T_725 ? issue_slots_10_uop_is_unique : _GEN_5775; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_sys_pc2epc = slots_10_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5974 = _T_725 ? issue_slots_10_uop_is_sys_pc2epc : _GEN_5776; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_uses_stq = slots_10_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5975 = _T_725 ? issue_slots_10_uop_uses_stq : _GEN_5777; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_uses_ldq = slots_10_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5976 = _T_725 ? issue_slots_10_uop_uses_ldq : _GEN_5778; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_amo = slots_10_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5977 = _T_725 ? issue_slots_10_uop_is_amo : _GEN_5779; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_fencei = slots_10_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5978 = _T_725 ? issue_slots_10_uop_is_fencei : _GEN_5780; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_fence = slots_10_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5979 = _T_725 ? issue_slots_10_uop_is_fence : _GEN_5781; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_mem_signed = slots_10_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5980 = _T_725 ? issue_slots_10_uop_mem_signed : _GEN_5782; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_mem_size = slots_10_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5981 = _T_725 ? issue_slots_10_uop_mem_size : _GEN_5783; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_mem_cmd = slots_10_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5982 = _T_725 ? issue_slots_10_uop_mem_cmd : _GEN_5784; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_bypassable = slots_10_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5983 = _T_725 ? issue_slots_10_uop_bypassable : _GEN_5785; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_10_uop_exc_cause = slots_10_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_5984 = _T_725 ? issue_slots_10_uop_exc_cause : _GEN_5786; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_exception = slots_10_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5985 = _T_725 ? issue_slots_10_uop_exception : _GEN_5787; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_stale_pdst = slots_10_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5986 = _T_725 ? issue_slots_10_uop_stale_pdst : _GEN_5788; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ppred_busy = slots_10_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5987 = _T_725 ? issue_slots_10_uop_ppred_busy : _GEN_5789; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_prs3_busy = slots_10_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5988 = _T_725 ? issue_slots_10_uop_prs3_busy : _GEN_5790; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_prs2_busy = slots_10_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5989 = _T_725 ? issue_slots_10_uop_prs2_busy : _GEN_5791; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_prs1_busy = slots_10_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_5990 = _T_725 ? issue_slots_10_uop_prs1_busy : _GEN_5792; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_ppred = slots_10_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5991 = _T_725 ? issue_slots_10_uop_ppred : _GEN_5793; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_prs3 = slots_10_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5992 = _T_725 ? issue_slots_10_uop_prs3 : _GEN_5794; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_prs2 = slots_10_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5993 = _T_725 ? issue_slots_10_uop_prs2 : _GEN_5795; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_prs1 = slots_10_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5994 = _T_725 ? issue_slots_10_uop_prs1 : _GEN_5796; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_pdst = slots_10_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_5995 = _T_725 ? issue_slots_10_uop_pdst : _GEN_5797; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_rxq_idx = slots_10_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_5996 = _T_725 ? issue_slots_10_uop_rxq_idx : _GEN_5798; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_stq_idx = slots_10_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5997 = _T_725 ? issue_slots_10_uop_stq_idx : _GEN_5799; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_ldq_idx = slots_10_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_5998 = _T_725 ? issue_slots_10_uop_ldq_idx : _GEN_5800; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_rob_idx = slots_10_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_5999 = _T_725 ? issue_slots_10_uop_rob_idx : _GEN_5801; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_10_uop_csr_addr = slots_10_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6000 = _T_725 ? issue_slots_10_uop_csr_addr : _GEN_5802; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_10_uop_imm_packed = slots_10_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_6001 = _T_725 ? issue_slots_10_uop_imm_packed : _GEN_5803; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_taken = slots_10_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6002 = _T_725 ? issue_slots_10_uop_taken : _GEN_5804; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_pc_lob = slots_10_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6003 = _T_725 ? issue_slots_10_uop_pc_lob : _GEN_5805; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_edge_inst = slots_10_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6004 = _T_725 ? issue_slots_10_uop_edge_inst : _GEN_5806; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_ftq_idx = slots_10_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6005 = _T_725 ? issue_slots_10_uop_ftq_idx : _GEN_5807; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_br_tag = slots_10_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6006 = _T_725 ? issue_slots_10_uop_br_tag : _GEN_5808; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_10_uop_br_mask = slots_10_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6007 = _T_725 ? issue_slots_10_uop_br_mask : _GEN_5809; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_sfb = slots_10_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6008 = _T_725 ? issue_slots_10_uop_is_sfb : _GEN_5810; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_jal = slots_10_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6009 = _T_725 ? issue_slots_10_uop_is_jal : _GEN_5811; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_jalr = slots_10_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6010 = _T_725 ? issue_slots_10_uop_is_jalr : _GEN_5812; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_br = slots_10_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6011 = _T_725 ? issue_slots_10_uop_is_br : _GEN_5813; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_iw_p2_poisoned = slots_10_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6012 = _T_725 ? issue_slots_10_uop_iw_p2_poisoned : _GEN_5814; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_iw_p1_poisoned = slots_10_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6013 = _T_725 ? issue_slots_10_uop_iw_p1_poisoned : _GEN_5815; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_iw_state = slots_10_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6014 = _T_725 ? issue_slots_10_uop_iw_state : _GEN_5816; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_ctrl_op3_sel = slots_10_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6015 = _T_725 ? issue_slots_10_uop_ctrl_op3_sel : _GEN_5817; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_is_std = slots_10_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6016 = _T_725 ? issue_slots_10_uop_ctrl_is_std : _GEN_5818; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_is_sta = slots_10_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6017 = _T_725 ? issue_slots_10_uop_ctrl_is_sta : _GEN_5819; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_is_load = slots_10_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6018 = _T_725 ? issue_slots_10_uop_ctrl_is_load : _GEN_5820; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_ctrl_csr_cmd = slots_10_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6019 = _T_725 ? issue_slots_10_uop_ctrl_csr_cmd : _GEN_5821; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_fcn_dw = slots_10_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6020 = _T_725 ? issue_slots_10_uop_ctrl_fcn_dw : _GEN_5822; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_ctrl_op_fcn = slots_10_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6021 = _T_725 ? issue_slots_10_uop_ctrl_op_fcn : _GEN_5823; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_ctrl_imm_sel = slots_10_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6022 = _T_725 ? issue_slots_10_uop_ctrl_imm_sel : _GEN_5824; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_ctrl_op2_sel = slots_10_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6023 = _T_725 ? issue_slots_10_uop_ctrl_op2_sel : _GEN_5825; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_ctrl_op1_sel = slots_10_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6024 = _T_725 ? issue_slots_10_uop_ctrl_op1_sel : _GEN_5826; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_ctrl_br_type = slots_10_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6025 = _T_725 ? issue_slots_10_uop_ctrl_br_type : _GEN_5827; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6026 = _T_725 ? issue_slots_10_uop_fu_code : _GEN_5828; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_iq_type = slots_10_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6027 = _T_725 ? issue_slots_10_uop_iq_type : _GEN_5829; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_10_uop_debug_pc = slots_10_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_6028 = _T_725 ? issue_slots_10_uop_debug_pc : _GEN_5830; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_rvc = slots_10_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6029 = _T_725 ? issue_slots_10_uop_is_rvc : _GEN_5831; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_10_uop_debug_inst = slots_10_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6030 = _T_725 ? issue_slots_10_uop_debug_inst : _GEN_5832; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_10_uop_inst = slots_10_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6031 = _T_725 ? issue_slots_10_uop_inst : _GEN_5833; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_uopc = slots_10_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6032 = _T_725 ? issue_slots_10_uop_uopc : _GEN_5834; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_address_num = slots_10_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6033 = _T_725 ? issue_slots_10_uop_address_num : _GEN_5835; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_rob_inst_idx = slots_10_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6034 = _T_725 ? issue_slots_10_uop_rob_inst_idx : _GEN_5836; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_self_index = slots_10_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6035 = _T_725 ? issue_slots_10_uop_self_index : _GEN_5837; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_split_num = slots_10_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6036 = _T_725 ? issue_slots_10_uop_split_num : _GEN_5838; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_op2_sel = slots_10_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6037 = _T_725 ? issue_slots_10_uop_op2_sel : _GEN_5839; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_op1_sel = slots_10_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6038 = _T_725 ? issue_slots_10_uop_op1_sel : _GEN_5840; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_stale_pflag = slots_10_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6039 = _T_725 ? issue_slots_10_uop_stale_pflag : _GEN_5841; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_pflag_busy = slots_10_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6040 = _T_725 ? issue_slots_10_uop_pflag_busy : _GEN_5842; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_pwflag = slots_10_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6041 = _T_725 ? issue_slots_10_uop_pwflag : _GEN_5843; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_prflag = slots_10_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6042 = _T_725 ? issue_slots_10_uop_prflag : _GEN_5844; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_wflag = slots_10_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6043 = _T_725 ? issue_slots_10_uop_wflag : _GEN_5845; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_rflag = slots_10_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6044 = _T_725 ? issue_slots_10_uop_rflag : _GEN_5846; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_lrs3_rtype = slots_10_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6045 = _T_725 ? issue_slots_10_uop_lrs3_rtype : _GEN_5847; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_shift = slots_10_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6046 = _T_725 ? issue_slots_10_uop_shift : _GEN_5848; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_unicore = slots_10_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6047 = _T_725 ? issue_slots_10_uop_is_unicore : _GEN_5849; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_switch_off = slots_10_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6048 = _T_725 ? issue_slots_10_uop_switch_off : _GEN_5850; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_switch = slots_10_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6049 = _T_725 ? issue_slots_10_uop_switch : _GEN_5851; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6052 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_debug_tsrc : _GEN_5854
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6053 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_debug_fsrc : _GEN_5855
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6054 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_bp_xcpt_if : _GEN_5856; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6055 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_bp_debug_if : _GEN_5857; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6056 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_xcpt_ma_if : _GEN_5858; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6057 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_xcpt_ae_if : _GEN_5859; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6058 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_xcpt_pf_if : _GEN_5860; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6059 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_fp_single : _GEN_5861; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6060 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_fp_val : _GEN_5862; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6061 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_frs3_en : _GEN_5863; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6062 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_lrs2_rtype : _GEN_5864
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6063 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_lrs1_rtype : _GEN_5865
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6064 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_dst_rtype : _GEN_5866; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6065 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ldst_val : _GEN_5867; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6066 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_lrs3 : _GEN_5868; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6067 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_lrs2 : _GEN_5869; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6068 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_lrs1 : _GEN_5870; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6069 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ldst : _GEN_5871; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6070 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ldst_is_rs1 : _GEN_5872; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6071 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_flush_on_commit : _GEN_5873
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6072 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_unique : _GEN_5874; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6073 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_sys_pc2epc : _GEN_5875; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6074 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_uses_stq : _GEN_5876; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6075 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_uses_ldq : _GEN_5877; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6076 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_amo : _GEN_5878; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6077 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_fencei : _GEN_5879; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6078 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_fence : _GEN_5880; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6079 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_mem_signed : _GEN_5881; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6080 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_mem_size : _GEN_5882; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6081 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_mem_cmd : _GEN_5883; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6082 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_bypassable : _GEN_5884; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_6083 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_exc_cause : _GEN_5885
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6084 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_exception : _GEN_5886; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6085 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_stale_pdst : _GEN_5887
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6086 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ppred_busy : _GEN_5888; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6087 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_prs3_busy : _GEN_5889; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6088 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_prs2_busy : _GEN_5890; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6089 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_prs1_busy : _GEN_5891; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6090 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ppred : _GEN_5892; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6091 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_prs3 : _GEN_5893; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6092 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_prs2 : _GEN_5894; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6093 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_prs1 : _GEN_5895; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6094 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_pdst : _GEN_5896; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6095 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_rxq_idx : _GEN_5897; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6096 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_stq_idx : _GEN_5898; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6097 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ldq_idx : _GEN_5899; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6098 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_rob_idx : _GEN_5900; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6099 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_csr_addr : _GEN_5901; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_6100 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_imm_packed :
    _GEN_5902; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6101 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_taken : _GEN_5903; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6102 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_pc_lob : _GEN_5904; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6103 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_edge_inst : _GEN_5905; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6104 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ftq_idx : _GEN_5906; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6105 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_br_tag : _GEN_5907; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6106 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_br_mask : _GEN_5908; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6107 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_sfb : _GEN_5909; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6108 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_jal : _GEN_5910; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6109 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_jalr : _GEN_5911; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6110 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_br : _GEN_5912; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6111 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_iw_p2_poisoned : _GEN_5913; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6112 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_iw_p1_poisoned : _GEN_5914; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6113 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_iw_state : _GEN_5915; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6114 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_op3_sel :
    _GEN_5916; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6115 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_is_std : _GEN_5917; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6116 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_is_sta : _GEN_5918; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6117 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_is_load : _GEN_5919; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6118 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_csr_cmd :
    _GEN_5920; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6119 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_fcn_dw : _GEN_5921; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6120 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_op_fcn :
    _GEN_5922; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6121 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_imm_sel :
    _GEN_5923; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6122 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_op2_sel :
    _GEN_5924; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6123 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_op1_sel :
    _GEN_5925; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6124 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_ctrl_br_type :
    _GEN_5926; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6125 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_fu_code : _GEN_5927; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6126 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_iq_type : _GEN_5928; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_6127 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_debug_pc : _GEN_5929; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6128 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_rvc : _GEN_5930; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6129 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_debug_inst :
    _GEN_5931; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6130 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_inst : _GEN_5932; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6131 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_uopc : _GEN_5933; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6132 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_address_num :
    _GEN_5934; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6133 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_rob_inst_idx :
    _GEN_5935; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6134 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_self_index : _GEN_5936
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6135 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_split_num : _GEN_5937; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6136 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_op2_sel : _GEN_5938; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6137 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_op1_sel : _GEN_5939; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6138 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_stale_pflag :
    _GEN_5940; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6139 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_pflag_busy : _GEN_5941; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6140 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_pwflag : _GEN_5942; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6141 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_prflag : _GEN_5943; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6142 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_wflag : _GEN_5944; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6143 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_rflag : _GEN_5945; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6144 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_lrs3_rtype : _GEN_5946
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6145 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_shift : _GEN_5947; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6146 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_is_unicore : _GEN_5948; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6147 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_switch_off : _GEN_5949; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6148 = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 ? issue_slots_10_uop_switch : _GEN_5950; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_debug_tsrc = slots_11_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6151 = _T_755 ? issue_slots_11_uop_debug_tsrc : _GEN_5953; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_debug_fsrc = slots_11_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6152 = _T_755 ? issue_slots_11_uop_debug_fsrc : _GEN_5954; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_bp_xcpt_if = slots_11_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6153 = _T_755 ? issue_slots_11_uop_bp_xcpt_if : _GEN_5955; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_bp_debug_if = slots_11_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6154 = _T_755 ? issue_slots_11_uop_bp_debug_if : _GEN_5956; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_xcpt_ma_if = slots_11_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6155 = _T_755 ? issue_slots_11_uop_xcpt_ma_if : _GEN_5957; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_xcpt_ae_if = slots_11_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6156 = _T_755 ? issue_slots_11_uop_xcpt_ae_if : _GEN_5958; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_xcpt_pf_if = slots_11_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6157 = _T_755 ? issue_slots_11_uop_xcpt_pf_if : _GEN_5959; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_fp_single = slots_11_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6158 = _T_755 ? issue_slots_11_uop_fp_single : _GEN_5960; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_fp_val = slots_11_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6159 = _T_755 ? issue_slots_11_uop_fp_val : _GEN_5961; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_frs3_en = slots_11_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6160 = _T_755 ? issue_slots_11_uop_frs3_en : _GEN_5962; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_lrs2_rtype = slots_11_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6161 = _T_755 ? issue_slots_11_uop_lrs2_rtype : _GEN_5963; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_lrs1_rtype = slots_11_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6162 = _T_755 ? issue_slots_11_uop_lrs1_rtype : _GEN_5964; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_dst_rtype = slots_11_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6163 = _T_755 ? issue_slots_11_uop_dst_rtype : _GEN_5965; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ldst_val = slots_11_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6164 = _T_755 ? issue_slots_11_uop_ldst_val : _GEN_5966; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_lrs3 = slots_11_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6165 = _T_755 ? issue_slots_11_uop_lrs3 : _GEN_5967; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_lrs2 = slots_11_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6166 = _T_755 ? issue_slots_11_uop_lrs2 : _GEN_5968; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_lrs1 = slots_11_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6167 = _T_755 ? issue_slots_11_uop_lrs1 : _GEN_5969; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_ldst = slots_11_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6168 = _T_755 ? issue_slots_11_uop_ldst : _GEN_5970; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ldst_is_rs1 = slots_11_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6169 = _T_755 ? issue_slots_11_uop_ldst_is_rs1 : _GEN_5971; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_flush_on_commit = slots_11_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6170 = _T_755 ? issue_slots_11_uop_flush_on_commit : _GEN_5972; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_unique = slots_11_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6171 = _T_755 ? issue_slots_11_uop_is_unique : _GEN_5973; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_sys_pc2epc = slots_11_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6172 = _T_755 ? issue_slots_11_uop_is_sys_pc2epc : _GEN_5974; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_uses_stq = slots_11_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6173 = _T_755 ? issue_slots_11_uop_uses_stq : _GEN_5975; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_uses_ldq = slots_11_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6174 = _T_755 ? issue_slots_11_uop_uses_ldq : _GEN_5976; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_amo = slots_11_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6175 = _T_755 ? issue_slots_11_uop_is_amo : _GEN_5977; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_fencei = slots_11_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6176 = _T_755 ? issue_slots_11_uop_is_fencei : _GEN_5978; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_fence = slots_11_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6177 = _T_755 ? issue_slots_11_uop_is_fence : _GEN_5979; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_mem_signed = slots_11_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6178 = _T_755 ? issue_slots_11_uop_mem_signed : _GEN_5980; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_mem_size = slots_11_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6179 = _T_755 ? issue_slots_11_uop_mem_size : _GEN_5981; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_mem_cmd = slots_11_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6180 = _T_755 ? issue_slots_11_uop_mem_cmd : _GEN_5982; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_bypassable = slots_11_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6181 = _T_755 ? issue_slots_11_uop_bypassable : _GEN_5983; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_11_uop_exc_cause = slots_11_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_6182 = _T_755 ? issue_slots_11_uop_exc_cause : _GEN_5984; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_exception = slots_11_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6183 = _T_755 ? issue_slots_11_uop_exception : _GEN_5985; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_stale_pdst = slots_11_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6184 = _T_755 ? issue_slots_11_uop_stale_pdst : _GEN_5986; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ppred_busy = slots_11_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6185 = _T_755 ? issue_slots_11_uop_ppred_busy : _GEN_5987; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_prs3_busy = slots_11_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6186 = _T_755 ? issue_slots_11_uop_prs3_busy : _GEN_5988; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_prs2_busy = slots_11_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6187 = _T_755 ? issue_slots_11_uop_prs2_busy : _GEN_5989; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_prs1_busy = slots_11_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6188 = _T_755 ? issue_slots_11_uop_prs1_busy : _GEN_5990; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_ppred = slots_11_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6189 = _T_755 ? issue_slots_11_uop_ppred : _GEN_5991; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_prs3 = slots_11_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6190 = _T_755 ? issue_slots_11_uop_prs3 : _GEN_5992; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_prs2 = slots_11_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6191 = _T_755 ? issue_slots_11_uop_prs2 : _GEN_5993; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_prs1 = slots_11_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6192 = _T_755 ? issue_slots_11_uop_prs1 : _GEN_5994; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_pdst = slots_11_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6193 = _T_755 ? issue_slots_11_uop_pdst : _GEN_5995; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_rxq_idx = slots_11_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6194 = _T_755 ? issue_slots_11_uop_rxq_idx : _GEN_5996; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_stq_idx = slots_11_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6195 = _T_755 ? issue_slots_11_uop_stq_idx : _GEN_5997; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_ldq_idx = slots_11_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6196 = _T_755 ? issue_slots_11_uop_ldq_idx : _GEN_5998; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_rob_idx = slots_11_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6197 = _T_755 ? issue_slots_11_uop_rob_idx : _GEN_5999; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_11_uop_csr_addr = slots_11_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6198 = _T_755 ? issue_slots_11_uop_csr_addr : _GEN_6000; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_11_uop_imm_packed = slots_11_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_6199 = _T_755 ? issue_slots_11_uop_imm_packed : _GEN_6001; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_taken = slots_11_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6200 = _T_755 ? issue_slots_11_uop_taken : _GEN_6002; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_pc_lob = slots_11_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6201 = _T_755 ? issue_slots_11_uop_pc_lob : _GEN_6003; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_edge_inst = slots_11_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6202 = _T_755 ? issue_slots_11_uop_edge_inst : _GEN_6004; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_ftq_idx = slots_11_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6203 = _T_755 ? issue_slots_11_uop_ftq_idx : _GEN_6005; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_br_tag = slots_11_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6204 = _T_755 ? issue_slots_11_uop_br_tag : _GEN_6006; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_11_uop_br_mask = slots_11_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6205 = _T_755 ? issue_slots_11_uop_br_mask : _GEN_6007; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_sfb = slots_11_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6206 = _T_755 ? issue_slots_11_uop_is_sfb : _GEN_6008; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_jal = slots_11_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6207 = _T_755 ? issue_slots_11_uop_is_jal : _GEN_6009; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_jalr = slots_11_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6208 = _T_755 ? issue_slots_11_uop_is_jalr : _GEN_6010; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_br = slots_11_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6209 = _T_755 ? issue_slots_11_uop_is_br : _GEN_6011; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_iw_p2_poisoned = slots_11_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6210 = _T_755 ? issue_slots_11_uop_iw_p2_poisoned : _GEN_6012; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_iw_p1_poisoned = slots_11_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6211 = _T_755 ? issue_slots_11_uop_iw_p1_poisoned : _GEN_6013; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_iw_state = slots_11_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6212 = _T_755 ? issue_slots_11_uop_iw_state : _GEN_6014; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_ctrl_op3_sel = slots_11_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6213 = _T_755 ? issue_slots_11_uop_ctrl_op3_sel : _GEN_6015; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_is_std = slots_11_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6214 = _T_755 ? issue_slots_11_uop_ctrl_is_std : _GEN_6016; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_is_sta = slots_11_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6215 = _T_755 ? issue_slots_11_uop_ctrl_is_sta : _GEN_6017; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_is_load = slots_11_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6216 = _T_755 ? issue_slots_11_uop_ctrl_is_load : _GEN_6018; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_ctrl_csr_cmd = slots_11_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6217 = _T_755 ? issue_slots_11_uop_ctrl_csr_cmd : _GEN_6019; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_fcn_dw = slots_11_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6218 = _T_755 ? issue_slots_11_uop_ctrl_fcn_dw : _GEN_6020; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_ctrl_op_fcn = slots_11_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6219 = _T_755 ? issue_slots_11_uop_ctrl_op_fcn : _GEN_6021; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_ctrl_imm_sel = slots_11_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6220 = _T_755 ? issue_slots_11_uop_ctrl_imm_sel : _GEN_6022; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_ctrl_op2_sel = slots_11_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6221 = _T_755 ? issue_slots_11_uop_ctrl_op2_sel : _GEN_6023; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_ctrl_op1_sel = slots_11_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6222 = _T_755 ? issue_slots_11_uop_ctrl_op1_sel : _GEN_6024; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_ctrl_br_type = slots_11_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6223 = _T_755 ? issue_slots_11_uop_ctrl_br_type : _GEN_6025; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6224 = _T_755 ? issue_slots_11_uop_fu_code : _GEN_6026; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_iq_type = slots_11_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6225 = _T_755 ? issue_slots_11_uop_iq_type : _GEN_6027; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_11_uop_debug_pc = slots_11_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_6226 = _T_755 ? issue_slots_11_uop_debug_pc : _GEN_6028; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_rvc = slots_11_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6227 = _T_755 ? issue_slots_11_uop_is_rvc : _GEN_6029; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_11_uop_debug_inst = slots_11_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6228 = _T_755 ? issue_slots_11_uop_debug_inst : _GEN_6030; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_11_uop_inst = slots_11_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6229 = _T_755 ? issue_slots_11_uop_inst : _GEN_6031; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_uopc = slots_11_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6230 = _T_755 ? issue_slots_11_uop_uopc : _GEN_6032; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_address_num = slots_11_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6231 = _T_755 ? issue_slots_11_uop_address_num : _GEN_6033; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_rob_inst_idx = slots_11_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6232 = _T_755 ? issue_slots_11_uop_rob_inst_idx : _GEN_6034; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_self_index = slots_11_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6233 = _T_755 ? issue_slots_11_uop_self_index : _GEN_6035; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_split_num = slots_11_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6234 = _T_755 ? issue_slots_11_uop_split_num : _GEN_6036; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_op2_sel = slots_11_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6235 = _T_755 ? issue_slots_11_uop_op2_sel : _GEN_6037; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_op1_sel = slots_11_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6236 = _T_755 ? issue_slots_11_uop_op1_sel : _GEN_6038; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_stale_pflag = slots_11_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6237 = _T_755 ? issue_slots_11_uop_stale_pflag : _GEN_6039; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_pflag_busy = slots_11_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6238 = _T_755 ? issue_slots_11_uop_pflag_busy : _GEN_6040; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_pwflag = slots_11_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6239 = _T_755 ? issue_slots_11_uop_pwflag : _GEN_6041; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_prflag = slots_11_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6240 = _T_755 ? issue_slots_11_uop_prflag : _GEN_6042; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_wflag = slots_11_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6241 = _T_755 ? issue_slots_11_uop_wflag : _GEN_6043; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_rflag = slots_11_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6242 = _T_755 ? issue_slots_11_uop_rflag : _GEN_6044; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_lrs3_rtype = slots_11_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6243 = _T_755 ? issue_slots_11_uop_lrs3_rtype : _GEN_6045; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_shift = slots_11_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6244 = _T_755 ? issue_slots_11_uop_shift : _GEN_6046; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_unicore = slots_11_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6245 = _T_755 ? issue_slots_11_uop_is_unicore : _GEN_6047; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_switch_off = slots_11_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6246 = _T_755 ? issue_slots_11_uop_switch_off : _GEN_6048; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_switch = slots_11_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6247 = _T_755 ? issue_slots_11_uop_switch : _GEN_6049; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6250 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_debug_tsrc : _GEN_6052
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6251 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_debug_fsrc : _GEN_6053
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6252 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_bp_xcpt_if : _GEN_6054; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6253 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_bp_debug_if : _GEN_6055; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6254 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_xcpt_ma_if : _GEN_6056; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6255 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_xcpt_ae_if : _GEN_6057; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6256 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_xcpt_pf_if : _GEN_6058; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6257 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_fp_single : _GEN_6059; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6258 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_fp_val : _GEN_6060; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6259 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_frs3_en : _GEN_6061; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6260 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_lrs2_rtype : _GEN_6062
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6261 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_lrs1_rtype : _GEN_6063
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6262 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_dst_rtype : _GEN_6064; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6263 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ldst_val : _GEN_6065; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6264 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_lrs3 : _GEN_6066; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6265 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_lrs2 : _GEN_6067; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6266 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_lrs1 : _GEN_6068; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6267 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ldst : _GEN_6069; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6268 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ldst_is_rs1 : _GEN_6070; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6269 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_flush_on_commit : _GEN_6071
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6270 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_unique : _GEN_6072; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6271 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_sys_pc2epc : _GEN_6073; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6272 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_uses_stq : _GEN_6074; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6273 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_uses_ldq : _GEN_6075; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6274 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_amo : _GEN_6076; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6275 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_fencei : _GEN_6077; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6276 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_fence : _GEN_6078; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6277 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_mem_signed : _GEN_6079; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6278 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_mem_size : _GEN_6080; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6279 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_mem_cmd : _GEN_6081; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6280 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_bypassable : _GEN_6082; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_6281 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_exc_cause : _GEN_6083
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6282 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_exception : _GEN_6084; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6283 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_stale_pdst : _GEN_6085
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6284 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ppred_busy : _GEN_6086; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6285 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_prs3_busy : _GEN_6087; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6286 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_prs2_busy : _GEN_6088; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6287 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_prs1_busy : _GEN_6089; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6288 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ppred : _GEN_6090; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6289 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_prs3 : _GEN_6091; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6290 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_prs2 : _GEN_6092; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6291 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_prs1 : _GEN_6093; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6292 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_pdst : _GEN_6094; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6293 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_rxq_idx : _GEN_6095; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6294 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_stq_idx : _GEN_6096; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6295 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ldq_idx : _GEN_6097; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6296 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_rob_idx : _GEN_6098; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6297 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_csr_addr : _GEN_6099; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_6298 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_imm_packed :
    _GEN_6100; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6299 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_taken : _GEN_6101; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6300 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_pc_lob : _GEN_6102; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6301 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_edge_inst : _GEN_6103; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6302 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ftq_idx : _GEN_6104; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6303 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_br_tag : _GEN_6105; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6304 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_br_mask : _GEN_6106; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6305 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_sfb : _GEN_6107; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6306 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_jal : _GEN_6108; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6307 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_jalr : _GEN_6109; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6308 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_br : _GEN_6110; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6309 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_iw_p2_poisoned : _GEN_6111; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6310 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_iw_p1_poisoned : _GEN_6112; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6311 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_iw_state : _GEN_6113; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6312 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_op3_sel :
    _GEN_6114; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6313 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_is_std : _GEN_6115; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6314 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_is_sta : _GEN_6116; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6315 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_is_load : _GEN_6117; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6316 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_csr_cmd :
    _GEN_6118; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6317 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_fcn_dw : _GEN_6119; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6318 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_op_fcn :
    _GEN_6120; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6319 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_imm_sel :
    _GEN_6121; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6320 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_op2_sel :
    _GEN_6122; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6321 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_op1_sel :
    _GEN_6123; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6322 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_ctrl_br_type :
    _GEN_6124; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6323 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_fu_code : _GEN_6125; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6324 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_iq_type : _GEN_6126; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_6325 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_debug_pc : _GEN_6127; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6326 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_rvc : _GEN_6128; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6327 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_debug_inst :
    _GEN_6129; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6328 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_inst : _GEN_6130; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6329 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_uopc : _GEN_6131; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6330 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_address_num :
    _GEN_6132; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6331 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_rob_inst_idx :
    _GEN_6133; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6332 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_self_index : _GEN_6134
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6333 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_split_num : _GEN_6135; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6334 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_op2_sel : _GEN_6136; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6335 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_op1_sel : _GEN_6137; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6336 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_stale_pflag :
    _GEN_6138; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6337 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_pflag_busy : _GEN_6139; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6338 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_pwflag : _GEN_6140; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6339 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_prflag : _GEN_6141; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6340 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_wflag : _GEN_6142; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6341 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_rflag : _GEN_6143; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6342 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_lrs3_rtype : _GEN_6144
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6343 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_shift : _GEN_6145; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6344 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_is_unicore : _GEN_6146; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6345 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_switch_off : _GEN_6147; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6346 = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 ? issue_slots_11_uop_switch : _GEN_6148; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_debug_tsrc = slots_12_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6349 = _T_785 ? issue_slots_12_uop_debug_tsrc : _GEN_6151; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_debug_fsrc = slots_12_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6350 = _T_785 ? issue_slots_12_uop_debug_fsrc : _GEN_6152; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_bp_xcpt_if = slots_12_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6351 = _T_785 ? issue_slots_12_uop_bp_xcpt_if : _GEN_6153; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_bp_debug_if = slots_12_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6352 = _T_785 ? issue_slots_12_uop_bp_debug_if : _GEN_6154; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_xcpt_ma_if = slots_12_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6353 = _T_785 ? issue_slots_12_uop_xcpt_ma_if : _GEN_6155; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_xcpt_ae_if = slots_12_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6354 = _T_785 ? issue_slots_12_uop_xcpt_ae_if : _GEN_6156; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_xcpt_pf_if = slots_12_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6355 = _T_785 ? issue_slots_12_uop_xcpt_pf_if : _GEN_6157; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_fp_single = slots_12_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6356 = _T_785 ? issue_slots_12_uop_fp_single : _GEN_6158; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_fp_val = slots_12_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6357 = _T_785 ? issue_slots_12_uop_fp_val : _GEN_6159; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_frs3_en = slots_12_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6358 = _T_785 ? issue_slots_12_uop_frs3_en : _GEN_6160; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_lrs2_rtype = slots_12_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6359 = _T_785 ? issue_slots_12_uop_lrs2_rtype : _GEN_6161; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_lrs1_rtype = slots_12_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6360 = _T_785 ? issue_slots_12_uop_lrs1_rtype : _GEN_6162; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_dst_rtype = slots_12_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6361 = _T_785 ? issue_slots_12_uop_dst_rtype : _GEN_6163; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ldst_val = slots_12_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6362 = _T_785 ? issue_slots_12_uop_ldst_val : _GEN_6164; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_lrs3 = slots_12_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6363 = _T_785 ? issue_slots_12_uop_lrs3 : _GEN_6165; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_lrs2 = slots_12_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6364 = _T_785 ? issue_slots_12_uop_lrs2 : _GEN_6166; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_lrs1 = slots_12_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6365 = _T_785 ? issue_slots_12_uop_lrs1 : _GEN_6167; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_ldst = slots_12_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6366 = _T_785 ? issue_slots_12_uop_ldst : _GEN_6168; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ldst_is_rs1 = slots_12_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6367 = _T_785 ? issue_slots_12_uop_ldst_is_rs1 : _GEN_6169; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_flush_on_commit = slots_12_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6368 = _T_785 ? issue_slots_12_uop_flush_on_commit : _GEN_6170; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_unique = slots_12_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6369 = _T_785 ? issue_slots_12_uop_is_unique : _GEN_6171; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_sys_pc2epc = slots_12_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6370 = _T_785 ? issue_slots_12_uop_is_sys_pc2epc : _GEN_6172; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_uses_stq = slots_12_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6371 = _T_785 ? issue_slots_12_uop_uses_stq : _GEN_6173; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_uses_ldq = slots_12_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6372 = _T_785 ? issue_slots_12_uop_uses_ldq : _GEN_6174; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_amo = slots_12_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6373 = _T_785 ? issue_slots_12_uop_is_amo : _GEN_6175; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_fencei = slots_12_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6374 = _T_785 ? issue_slots_12_uop_is_fencei : _GEN_6176; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_fence = slots_12_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6375 = _T_785 ? issue_slots_12_uop_is_fence : _GEN_6177; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_mem_signed = slots_12_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6376 = _T_785 ? issue_slots_12_uop_mem_signed : _GEN_6178; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_mem_size = slots_12_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6377 = _T_785 ? issue_slots_12_uop_mem_size : _GEN_6179; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_mem_cmd = slots_12_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6378 = _T_785 ? issue_slots_12_uop_mem_cmd : _GEN_6180; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_bypassable = slots_12_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6379 = _T_785 ? issue_slots_12_uop_bypassable : _GEN_6181; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_12_uop_exc_cause = slots_12_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_6380 = _T_785 ? issue_slots_12_uop_exc_cause : _GEN_6182; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_exception = slots_12_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6381 = _T_785 ? issue_slots_12_uop_exception : _GEN_6183; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_stale_pdst = slots_12_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6382 = _T_785 ? issue_slots_12_uop_stale_pdst : _GEN_6184; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ppred_busy = slots_12_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6383 = _T_785 ? issue_slots_12_uop_ppred_busy : _GEN_6185; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_prs3_busy = slots_12_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6384 = _T_785 ? issue_slots_12_uop_prs3_busy : _GEN_6186; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_prs2_busy = slots_12_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6385 = _T_785 ? issue_slots_12_uop_prs2_busy : _GEN_6187; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_prs1_busy = slots_12_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6386 = _T_785 ? issue_slots_12_uop_prs1_busy : _GEN_6188; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_ppred = slots_12_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6387 = _T_785 ? issue_slots_12_uop_ppred : _GEN_6189; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_prs3 = slots_12_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6388 = _T_785 ? issue_slots_12_uop_prs3 : _GEN_6190; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_prs2 = slots_12_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6389 = _T_785 ? issue_slots_12_uop_prs2 : _GEN_6191; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_prs1 = slots_12_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6390 = _T_785 ? issue_slots_12_uop_prs1 : _GEN_6192; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_pdst = slots_12_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6391 = _T_785 ? issue_slots_12_uop_pdst : _GEN_6193; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_rxq_idx = slots_12_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6392 = _T_785 ? issue_slots_12_uop_rxq_idx : _GEN_6194; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_stq_idx = slots_12_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6393 = _T_785 ? issue_slots_12_uop_stq_idx : _GEN_6195; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_ldq_idx = slots_12_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6394 = _T_785 ? issue_slots_12_uop_ldq_idx : _GEN_6196; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_rob_idx = slots_12_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6395 = _T_785 ? issue_slots_12_uop_rob_idx : _GEN_6197; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_12_uop_csr_addr = slots_12_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6396 = _T_785 ? issue_slots_12_uop_csr_addr : _GEN_6198; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_12_uop_imm_packed = slots_12_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_6397 = _T_785 ? issue_slots_12_uop_imm_packed : _GEN_6199; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_taken = slots_12_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6398 = _T_785 ? issue_slots_12_uop_taken : _GEN_6200; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_pc_lob = slots_12_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6399 = _T_785 ? issue_slots_12_uop_pc_lob : _GEN_6201; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_edge_inst = slots_12_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6400 = _T_785 ? issue_slots_12_uop_edge_inst : _GEN_6202; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_ftq_idx = slots_12_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6401 = _T_785 ? issue_slots_12_uop_ftq_idx : _GEN_6203; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_br_tag = slots_12_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6402 = _T_785 ? issue_slots_12_uop_br_tag : _GEN_6204; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_12_uop_br_mask = slots_12_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6403 = _T_785 ? issue_slots_12_uop_br_mask : _GEN_6205; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_sfb = slots_12_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6404 = _T_785 ? issue_slots_12_uop_is_sfb : _GEN_6206; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_jal = slots_12_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6405 = _T_785 ? issue_slots_12_uop_is_jal : _GEN_6207; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_jalr = slots_12_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6406 = _T_785 ? issue_slots_12_uop_is_jalr : _GEN_6208; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_br = slots_12_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6407 = _T_785 ? issue_slots_12_uop_is_br : _GEN_6209; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_iw_p2_poisoned = slots_12_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6408 = _T_785 ? issue_slots_12_uop_iw_p2_poisoned : _GEN_6210; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_iw_p1_poisoned = slots_12_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6409 = _T_785 ? issue_slots_12_uop_iw_p1_poisoned : _GEN_6211; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_iw_state = slots_12_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6410 = _T_785 ? issue_slots_12_uop_iw_state : _GEN_6212; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_ctrl_op3_sel = slots_12_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6411 = _T_785 ? issue_slots_12_uop_ctrl_op3_sel : _GEN_6213; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_is_std = slots_12_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6412 = _T_785 ? issue_slots_12_uop_ctrl_is_std : _GEN_6214; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_is_sta = slots_12_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6413 = _T_785 ? issue_slots_12_uop_ctrl_is_sta : _GEN_6215; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_is_load = slots_12_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6414 = _T_785 ? issue_slots_12_uop_ctrl_is_load : _GEN_6216; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_ctrl_csr_cmd = slots_12_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6415 = _T_785 ? issue_slots_12_uop_ctrl_csr_cmd : _GEN_6217; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_fcn_dw = slots_12_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6416 = _T_785 ? issue_slots_12_uop_ctrl_fcn_dw : _GEN_6218; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_ctrl_op_fcn = slots_12_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6417 = _T_785 ? issue_slots_12_uop_ctrl_op_fcn : _GEN_6219; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_ctrl_imm_sel = slots_12_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6418 = _T_785 ? issue_slots_12_uop_ctrl_imm_sel : _GEN_6220; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_ctrl_op2_sel = slots_12_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6419 = _T_785 ? issue_slots_12_uop_ctrl_op2_sel : _GEN_6221; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_ctrl_op1_sel = slots_12_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6420 = _T_785 ? issue_slots_12_uop_ctrl_op1_sel : _GEN_6222; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_ctrl_br_type = slots_12_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6421 = _T_785 ? issue_slots_12_uop_ctrl_br_type : _GEN_6223; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6422 = _T_785 ? issue_slots_12_uop_fu_code : _GEN_6224; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_iq_type = slots_12_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6423 = _T_785 ? issue_slots_12_uop_iq_type : _GEN_6225; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_12_uop_debug_pc = slots_12_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_6424 = _T_785 ? issue_slots_12_uop_debug_pc : _GEN_6226; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_rvc = slots_12_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6425 = _T_785 ? issue_slots_12_uop_is_rvc : _GEN_6227; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_12_uop_debug_inst = slots_12_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6426 = _T_785 ? issue_slots_12_uop_debug_inst : _GEN_6228; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_12_uop_inst = slots_12_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6427 = _T_785 ? issue_slots_12_uop_inst : _GEN_6229; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_uopc = slots_12_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6428 = _T_785 ? issue_slots_12_uop_uopc : _GEN_6230; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_address_num = slots_12_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6429 = _T_785 ? issue_slots_12_uop_address_num : _GEN_6231; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_rob_inst_idx = slots_12_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6430 = _T_785 ? issue_slots_12_uop_rob_inst_idx : _GEN_6232; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_self_index = slots_12_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6431 = _T_785 ? issue_slots_12_uop_self_index : _GEN_6233; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_split_num = slots_12_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6432 = _T_785 ? issue_slots_12_uop_split_num : _GEN_6234; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_op2_sel = slots_12_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6433 = _T_785 ? issue_slots_12_uop_op2_sel : _GEN_6235; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_op1_sel = slots_12_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6434 = _T_785 ? issue_slots_12_uop_op1_sel : _GEN_6236; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_stale_pflag = slots_12_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6435 = _T_785 ? issue_slots_12_uop_stale_pflag : _GEN_6237; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_pflag_busy = slots_12_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6436 = _T_785 ? issue_slots_12_uop_pflag_busy : _GEN_6238; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_pwflag = slots_12_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6437 = _T_785 ? issue_slots_12_uop_pwflag : _GEN_6239; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_prflag = slots_12_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6438 = _T_785 ? issue_slots_12_uop_prflag : _GEN_6240; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_wflag = slots_12_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6439 = _T_785 ? issue_slots_12_uop_wflag : _GEN_6241; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_rflag = slots_12_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6440 = _T_785 ? issue_slots_12_uop_rflag : _GEN_6242; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_lrs3_rtype = slots_12_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6441 = _T_785 ? issue_slots_12_uop_lrs3_rtype : _GEN_6243; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_shift = slots_12_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6442 = _T_785 ? issue_slots_12_uop_shift : _GEN_6244; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_unicore = slots_12_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6443 = _T_785 ? issue_slots_12_uop_is_unicore : _GEN_6245; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_switch_off = slots_12_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6444 = _T_785 ? issue_slots_12_uop_switch_off : _GEN_6246; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_switch = slots_12_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6445 = _T_785 ? issue_slots_12_uop_switch : _GEN_6247; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6448 = _T_796 & ~_T_767 ? issue_slots_12_uop_debug_tsrc : _GEN_6250; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6449 = _T_796 & ~_T_767 ? issue_slots_12_uop_debug_fsrc : _GEN_6251; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6450 = _T_796 & ~_T_767 ? issue_slots_12_uop_bp_xcpt_if : _GEN_6252; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6451 = _T_796 & ~_T_767 ? issue_slots_12_uop_bp_debug_if : _GEN_6253; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6452 = _T_796 & ~_T_767 ? issue_slots_12_uop_xcpt_ma_if : _GEN_6254; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6453 = _T_796 & ~_T_767 ? issue_slots_12_uop_xcpt_ae_if : _GEN_6255; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6454 = _T_796 & ~_T_767 ? issue_slots_12_uop_xcpt_pf_if : _GEN_6256; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6455 = _T_796 & ~_T_767 ? issue_slots_12_uop_fp_single : _GEN_6257; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6456 = _T_796 & ~_T_767 ? issue_slots_12_uop_fp_val : _GEN_6258; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6457 = _T_796 & ~_T_767 ? issue_slots_12_uop_frs3_en : _GEN_6259; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6458 = _T_796 & ~_T_767 ? issue_slots_12_uop_lrs2_rtype : _GEN_6260; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6459 = _T_796 & ~_T_767 ? issue_slots_12_uop_lrs1_rtype : _GEN_6261; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6460 = _T_796 & ~_T_767 ? issue_slots_12_uop_dst_rtype : _GEN_6262; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6461 = _T_796 & ~_T_767 ? issue_slots_12_uop_ldst_val : _GEN_6263; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6462 = _T_796 & ~_T_767 ? issue_slots_12_uop_lrs3 : _GEN_6264; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6463 = _T_796 & ~_T_767 ? issue_slots_12_uop_lrs2 : _GEN_6265; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6464 = _T_796 & ~_T_767 ? issue_slots_12_uop_lrs1 : _GEN_6266; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6465 = _T_796 & ~_T_767 ? issue_slots_12_uop_ldst : _GEN_6267; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6466 = _T_796 & ~_T_767 ? issue_slots_12_uop_ldst_is_rs1 : _GEN_6268; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6467 = _T_796 & ~_T_767 ? issue_slots_12_uop_flush_on_commit : _GEN_6269; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6468 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_unique : _GEN_6270; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6469 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_sys_pc2epc : _GEN_6271; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6470 = _T_796 & ~_T_767 ? issue_slots_12_uop_uses_stq : _GEN_6272; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6471 = _T_796 & ~_T_767 ? issue_slots_12_uop_uses_ldq : _GEN_6273; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6472 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_amo : _GEN_6274; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6473 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_fencei : _GEN_6275; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6474 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_fence : _GEN_6276; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6475 = _T_796 & ~_T_767 ? issue_slots_12_uop_mem_signed : _GEN_6277; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6476 = _T_796 & ~_T_767 ? issue_slots_12_uop_mem_size : _GEN_6278; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6477 = _T_796 & ~_T_767 ? issue_slots_12_uop_mem_cmd : _GEN_6279; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6478 = _T_796 & ~_T_767 ? issue_slots_12_uop_bypassable : _GEN_6280; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_6479 = _T_796 & ~_T_767 ? issue_slots_12_uop_exc_cause : _GEN_6281; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6480 = _T_796 & ~_T_767 ? issue_slots_12_uop_exception : _GEN_6282; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6481 = _T_796 & ~_T_767 ? issue_slots_12_uop_stale_pdst : _GEN_6283; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6482 = _T_796 & ~_T_767 ? issue_slots_12_uop_ppred_busy : _GEN_6284; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6483 = _T_796 & ~_T_767 ? issue_slots_12_uop_prs3_busy : _GEN_6285; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6484 = _T_796 & ~_T_767 ? issue_slots_12_uop_prs2_busy : _GEN_6286; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6485 = _T_796 & ~_T_767 ? issue_slots_12_uop_prs1_busy : _GEN_6287; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6486 = _T_796 & ~_T_767 ? issue_slots_12_uop_ppred : _GEN_6288; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6487 = _T_796 & ~_T_767 ? issue_slots_12_uop_prs3 : _GEN_6289; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6488 = _T_796 & ~_T_767 ? issue_slots_12_uop_prs2 : _GEN_6290; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6489 = _T_796 & ~_T_767 ? issue_slots_12_uop_prs1 : _GEN_6291; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6490 = _T_796 & ~_T_767 ? issue_slots_12_uop_pdst : _GEN_6292; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6491 = _T_796 & ~_T_767 ? issue_slots_12_uop_rxq_idx : _GEN_6293; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6492 = _T_796 & ~_T_767 ? issue_slots_12_uop_stq_idx : _GEN_6294; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6493 = _T_796 & ~_T_767 ? issue_slots_12_uop_ldq_idx : _GEN_6295; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6494 = _T_796 & ~_T_767 ? issue_slots_12_uop_rob_idx : _GEN_6296; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6495 = _T_796 & ~_T_767 ? issue_slots_12_uop_csr_addr : _GEN_6297; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_6496 = _T_796 & ~_T_767 ? issue_slots_12_uop_imm_packed : _GEN_6298; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6497 = _T_796 & ~_T_767 ? issue_slots_12_uop_taken : _GEN_6299; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6498 = _T_796 & ~_T_767 ? issue_slots_12_uop_pc_lob : _GEN_6300; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6499 = _T_796 & ~_T_767 ? issue_slots_12_uop_edge_inst : _GEN_6301; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6500 = _T_796 & ~_T_767 ? issue_slots_12_uop_ftq_idx : _GEN_6302; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6501 = _T_796 & ~_T_767 ? issue_slots_12_uop_br_tag : _GEN_6303; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6502 = _T_796 & ~_T_767 ? issue_slots_12_uop_br_mask : _GEN_6304; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6503 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_sfb : _GEN_6305; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6504 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_jal : _GEN_6306; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6505 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_jalr : _GEN_6307; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6506 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_br : _GEN_6308; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6507 = _T_796 & ~_T_767 ? issue_slots_12_uop_iw_p2_poisoned : _GEN_6309; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6508 = _T_796 & ~_T_767 ? issue_slots_12_uop_iw_p1_poisoned : _GEN_6310; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6509 = _T_796 & ~_T_767 ? issue_slots_12_uop_iw_state : _GEN_6311; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6510 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_op3_sel : _GEN_6312; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6511 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_is_std : _GEN_6313; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6512 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_is_sta : _GEN_6314; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6513 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_is_load : _GEN_6315; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6514 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_csr_cmd : _GEN_6316; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6515 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_fcn_dw : _GEN_6317; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6516 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_op_fcn : _GEN_6318; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6517 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_imm_sel : _GEN_6319; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6518 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_op2_sel : _GEN_6320; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6519 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_op1_sel : _GEN_6321; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6520 = _T_796 & ~_T_767 ? issue_slots_12_uop_ctrl_br_type : _GEN_6322; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6521 = _T_796 & ~_T_767 ? issue_slots_12_uop_fu_code : _GEN_6323; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6522 = _T_796 & ~_T_767 ? issue_slots_12_uop_iq_type : _GEN_6324; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_6523 = _T_796 & ~_T_767 ? issue_slots_12_uop_debug_pc : _GEN_6325; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6524 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_rvc : _GEN_6326; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6525 = _T_796 & ~_T_767 ? issue_slots_12_uop_debug_inst : _GEN_6327; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6526 = _T_796 & ~_T_767 ? issue_slots_12_uop_inst : _GEN_6328; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6527 = _T_796 & ~_T_767 ? issue_slots_12_uop_uopc : _GEN_6329; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6528 = _T_796 & ~_T_767 ? issue_slots_12_uop_address_num : _GEN_6330; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6529 = _T_796 & ~_T_767 ? issue_slots_12_uop_rob_inst_idx : _GEN_6331; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6530 = _T_796 & ~_T_767 ? issue_slots_12_uop_self_index : _GEN_6332; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6531 = _T_796 & ~_T_767 ? issue_slots_12_uop_split_num : _GEN_6333; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6532 = _T_796 & ~_T_767 ? issue_slots_12_uop_op2_sel : _GEN_6334; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6533 = _T_796 & ~_T_767 ? issue_slots_12_uop_op1_sel : _GEN_6335; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6534 = _T_796 & ~_T_767 ? issue_slots_12_uop_stale_pflag : _GEN_6336; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6535 = _T_796 & ~_T_767 ? issue_slots_12_uop_pflag_busy : _GEN_6337; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6536 = _T_796 & ~_T_767 ? issue_slots_12_uop_pwflag : _GEN_6338; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6537 = _T_796 & ~_T_767 ? issue_slots_12_uop_prflag : _GEN_6339; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6538 = _T_796 & ~_T_767 ? issue_slots_12_uop_wflag : _GEN_6340; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6539 = _T_796 & ~_T_767 ? issue_slots_12_uop_rflag : _GEN_6341; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6540 = _T_796 & ~_T_767 ? issue_slots_12_uop_lrs3_rtype : _GEN_6342; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6541 = _T_796 & ~_T_767 ? issue_slots_12_uop_shift : _GEN_6343; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6542 = _T_796 & ~_T_767 ? issue_slots_12_uop_is_unicore : _GEN_6344; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6543 = _T_796 & ~_T_767 ? issue_slots_12_uop_switch_off : _GEN_6345; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6544 = _T_796 & ~_T_767 ? issue_slots_12_uop_switch : _GEN_6346; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_debug_tsrc = slots_13_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6547 = _T_815 ? issue_slots_13_uop_debug_tsrc : _GEN_6349; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_debug_fsrc = slots_13_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6548 = _T_815 ? issue_slots_13_uop_debug_fsrc : _GEN_6350; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_bp_xcpt_if = slots_13_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6549 = _T_815 ? issue_slots_13_uop_bp_xcpt_if : _GEN_6351; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_bp_debug_if = slots_13_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6550 = _T_815 ? issue_slots_13_uop_bp_debug_if : _GEN_6352; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_xcpt_ma_if = slots_13_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6551 = _T_815 ? issue_slots_13_uop_xcpt_ma_if : _GEN_6353; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_xcpt_ae_if = slots_13_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6552 = _T_815 ? issue_slots_13_uop_xcpt_ae_if : _GEN_6354; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_xcpt_pf_if = slots_13_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6553 = _T_815 ? issue_slots_13_uop_xcpt_pf_if : _GEN_6355; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_fp_single = slots_13_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6554 = _T_815 ? issue_slots_13_uop_fp_single : _GEN_6356; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_fp_val = slots_13_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6555 = _T_815 ? issue_slots_13_uop_fp_val : _GEN_6357; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_frs3_en = slots_13_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6556 = _T_815 ? issue_slots_13_uop_frs3_en : _GEN_6358; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_lrs2_rtype = slots_13_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6557 = _T_815 ? issue_slots_13_uop_lrs2_rtype : _GEN_6359; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_lrs1_rtype = slots_13_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6558 = _T_815 ? issue_slots_13_uop_lrs1_rtype : _GEN_6360; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_dst_rtype = slots_13_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6559 = _T_815 ? issue_slots_13_uop_dst_rtype : _GEN_6361; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ldst_val = slots_13_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6560 = _T_815 ? issue_slots_13_uop_ldst_val : _GEN_6362; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_lrs3 = slots_13_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6561 = _T_815 ? issue_slots_13_uop_lrs3 : _GEN_6363; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_lrs2 = slots_13_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6562 = _T_815 ? issue_slots_13_uop_lrs2 : _GEN_6364; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_lrs1 = slots_13_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6563 = _T_815 ? issue_slots_13_uop_lrs1 : _GEN_6365; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_ldst = slots_13_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6564 = _T_815 ? issue_slots_13_uop_ldst : _GEN_6366; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ldst_is_rs1 = slots_13_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6565 = _T_815 ? issue_slots_13_uop_ldst_is_rs1 : _GEN_6367; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_flush_on_commit = slots_13_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6566 = _T_815 ? issue_slots_13_uop_flush_on_commit : _GEN_6368; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_unique = slots_13_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6567 = _T_815 ? issue_slots_13_uop_is_unique : _GEN_6369; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_sys_pc2epc = slots_13_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6568 = _T_815 ? issue_slots_13_uop_is_sys_pc2epc : _GEN_6370; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_uses_stq = slots_13_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6569 = _T_815 ? issue_slots_13_uop_uses_stq : _GEN_6371; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_uses_ldq = slots_13_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6570 = _T_815 ? issue_slots_13_uop_uses_ldq : _GEN_6372; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_amo = slots_13_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6571 = _T_815 ? issue_slots_13_uop_is_amo : _GEN_6373; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_fencei = slots_13_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6572 = _T_815 ? issue_slots_13_uop_is_fencei : _GEN_6374; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_fence = slots_13_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6573 = _T_815 ? issue_slots_13_uop_is_fence : _GEN_6375; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_mem_signed = slots_13_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6574 = _T_815 ? issue_slots_13_uop_mem_signed : _GEN_6376; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_mem_size = slots_13_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6575 = _T_815 ? issue_slots_13_uop_mem_size : _GEN_6377; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_mem_cmd = slots_13_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6576 = _T_815 ? issue_slots_13_uop_mem_cmd : _GEN_6378; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_bypassable = slots_13_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6577 = _T_815 ? issue_slots_13_uop_bypassable : _GEN_6379; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_13_uop_exc_cause = slots_13_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_6578 = _T_815 ? issue_slots_13_uop_exc_cause : _GEN_6380; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_exception = slots_13_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6579 = _T_815 ? issue_slots_13_uop_exception : _GEN_6381; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_stale_pdst = slots_13_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6580 = _T_815 ? issue_slots_13_uop_stale_pdst : _GEN_6382; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ppred_busy = slots_13_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6581 = _T_815 ? issue_slots_13_uop_ppred_busy : _GEN_6383; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_prs3_busy = slots_13_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6582 = _T_815 ? issue_slots_13_uop_prs3_busy : _GEN_6384; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_prs2_busy = slots_13_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6583 = _T_815 ? issue_slots_13_uop_prs2_busy : _GEN_6385; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_prs1_busy = slots_13_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6584 = _T_815 ? issue_slots_13_uop_prs1_busy : _GEN_6386; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_ppred = slots_13_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6585 = _T_815 ? issue_slots_13_uop_ppred : _GEN_6387; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_prs3 = slots_13_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6586 = _T_815 ? issue_slots_13_uop_prs3 : _GEN_6388; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_prs2 = slots_13_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6587 = _T_815 ? issue_slots_13_uop_prs2 : _GEN_6389; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_prs1 = slots_13_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6588 = _T_815 ? issue_slots_13_uop_prs1 : _GEN_6390; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_pdst = slots_13_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6589 = _T_815 ? issue_slots_13_uop_pdst : _GEN_6391; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_rxq_idx = slots_13_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6590 = _T_815 ? issue_slots_13_uop_rxq_idx : _GEN_6392; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_stq_idx = slots_13_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6591 = _T_815 ? issue_slots_13_uop_stq_idx : _GEN_6393; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_ldq_idx = slots_13_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6592 = _T_815 ? issue_slots_13_uop_ldq_idx : _GEN_6394; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_rob_idx = slots_13_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6593 = _T_815 ? issue_slots_13_uop_rob_idx : _GEN_6395; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_13_uop_csr_addr = slots_13_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6594 = _T_815 ? issue_slots_13_uop_csr_addr : _GEN_6396; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_13_uop_imm_packed = slots_13_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_6595 = _T_815 ? issue_slots_13_uop_imm_packed : _GEN_6397; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_taken = slots_13_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6596 = _T_815 ? issue_slots_13_uop_taken : _GEN_6398; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_pc_lob = slots_13_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6597 = _T_815 ? issue_slots_13_uop_pc_lob : _GEN_6399; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_edge_inst = slots_13_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6598 = _T_815 ? issue_slots_13_uop_edge_inst : _GEN_6400; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_ftq_idx = slots_13_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6599 = _T_815 ? issue_slots_13_uop_ftq_idx : _GEN_6401; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_br_tag = slots_13_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6600 = _T_815 ? issue_slots_13_uop_br_tag : _GEN_6402; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_13_uop_br_mask = slots_13_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6601 = _T_815 ? issue_slots_13_uop_br_mask : _GEN_6403; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_sfb = slots_13_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6602 = _T_815 ? issue_slots_13_uop_is_sfb : _GEN_6404; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_jal = slots_13_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6603 = _T_815 ? issue_slots_13_uop_is_jal : _GEN_6405; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_jalr = slots_13_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6604 = _T_815 ? issue_slots_13_uop_is_jalr : _GEN_6406; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_br = slots_13_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6605 = _T_815 ? issue_slots_13_uop_is_br : _GEN_6407; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_iw_p2_poisoned = slots_13_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6606 = _T_815 ? issue_slots_13_uop_iw_p2_poisoned : _GEN_6408; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_iw_p1_poisoned = slots_13_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6607 = _T_815 ? issue_slots_13_uop_iw_p1_poisoned : _GEN_6409; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_iw_state = slots_13_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6608 = _T_815 ? issue_slots_13_uop_iw_state : _GEN_6410; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_ctrl_op3_sel = slots_13_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6609 = _T_815 ? issue_slots_13_uop_ctrl_op3_sel : _GEN_6411; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_is_std = slots_13_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6610 = _T_815 ? issue_slots_13_uop_ctrl_is_std : _GEN_6412; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_is_sta = slots_13_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6611 = _T_815 ? issue_slots_13_uop_ctrl_is_sta : _GEN_6413; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_is_load = slots_13_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6612 = _T_815 ? issue_slots_13_uop_ctrl_is_load : _GEN_6414; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_ctrl_csr_cmd = slots_13_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6613 = _T_815 ? issue_slots_13_uop_ctrl_csr_cmd : _GEN_6415; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_fcn_dw = slots_13_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6614 = _T_815 ? issue_slots_13_uop_ctrl_fcn_dw : _GEN_6416; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_ctrl_op_fcn = slots_13_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6615 = _T_815 ? issue_slots_13_uop_ctrl_op_fcn : _GEN_6417; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_ctrl_imm_sel = slots_13_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6616 = _T_815 ? issue_slots_13_uop_ctrl_imm_sel : _GEN_6418; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_ctrl_op2_sel = slots_13_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6617 = _T_815 ? issue_slots_13_uop_ctrl_op2_sel : _GEN_6419; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_ctrl_op1_sel = slots_13_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6618 = _T_815 ? issue_slots_13_uop_ctrl_op1_sel : _GEN_6420; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_ctrl_br_type = slots_13_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6619 = _T_815 ? issue_slots_13_uop_ctrl_br_type : _GEN_6421; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6620 = _T_815 ? issue_slots_13_uop_fu_code : _GEN_6422; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_iq_type = slots_13_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6621 = _T_815 ? issue_slots_13_uop_iq_type : _GEN_6423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_13_uop_debug_pc = slots_13_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_6622 = _T_815 ? issue_slots_13_uop_debug_pc : _GEN_6424; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_rvc = slots_13_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6623 = _T_815 ? issue_slots_13_uop_is_rvc : _GEN_6425; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_13_uop_debug_inst = slots_13_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6624 = _T_815 ? issue_slots_13_uop_debug_inst : _GEN_6426; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_13_uop_inst = slots_13_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6625 = _T_815 ? issue_slots_13_uop_inst : _GEN_6427; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_uopc = slots_13_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6626 = _T_815 ? issue_slots_13_uop_uopc : _GEN_6428; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_address_num = slots_13_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6627 = _T_815 ? issue_slots_13_uop_address_num : _GEN_6429; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_rob_inst_idx = slots_13_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6628 = _T_815 ? issue_slots_13_uop_rob_inst_idx : _GEN_6430; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_self_index = slots_13_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6629 = _T_815 ? issue_slots_13_uop_self_index : _GEN_6431; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_split_num = slots_13_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6630 = _T_815 ? issue_slots_13_uop_split_num : _GEN_6432; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_op2_sel = slots_13_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6631 = _T_815 ? issue_slots_13_uop_op2_sel : _GEN_6433; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_op1_sel = slots_13_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6632 = _T_815 ? issue_slots_13_uop_op1_sel : _GEN_6434; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_stale_pflag = slots_13_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6633 = _T_815 ? issue_slots_13_uop_stale_pflag : _GEN_6435; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_pflag_busy = slots_13_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6634 = _T_815 ? issue_slots_13_uop_pflag_busy : _GEN_6436; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_pwflag = slots_13_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6635 = _T_815 ? issue_slots_13_uop_pwflag : _GEN_6437; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_prflag = slots_13_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6636 = _T_815 ? issue_slots_13_uop_prflag : _GEN_6438; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_wflag = slots_13_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6637 = _T_815 ? issue_slots_13_uop_wflag : _GEN_6439; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_rflag = slots_13_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6638 = _T_815 ? issue_slots_13_uop_rflag : _GEN_6440; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_lrs3_rtype = slots_13_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6639 = _T_815 ? issue_slots_13_uop_lrs3_rtype : _GEN_6441; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_shift = slots_13_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6640 = _T_815 ? issue_slots_13_uop_shift : _GEN_6442; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_unicore = slots_13_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6641 = _T_815 ? issue_slots_13_uop_is_unicore : _GEN_6443; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_switch_off = slots_13_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6642 = _T_815 ? issue_slots_13_uop_switch_off : _GEN_6444; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_switch = slots_13_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6643 = _T_815 ? issue_slots_13_uop_switch : _GEN_6445; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6646 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_debug_tsrc : _GEN_6448
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6647 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_debug_fsrc : _GEN_6449
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6648 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_bp_xcpt_if : _GEN_6450; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6649 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_bp_debug_if : _GEN_6451; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6650 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_xcpt_ma_if : _GEN_6452; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6651 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_xcpt_ae_if : _GEN_6453; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6652 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_xcpt_pf_if : _GEN_6454; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6653 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_fp_single : _GEN_6455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6654 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_fp_val : _GEN_6456; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6655 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_frs3_en : _GEN_6457; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6656 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_lrs2_rtype : _GEN_6458
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6657 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_lrs1_rtype : _GEN_6459
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6658 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_dst_rtype : _GEN_6460; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6659 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ldst_val : _GEN_6461; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6660 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_lrs3 : _GEN_6462; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6661 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_lrs2 : _GEN_6463; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6662 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_lrs1 : _GEN_6464; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6663 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ldst : _GEN_6465; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6664 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ldst_is_rs1 : _GEN_6466; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6665 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_flush_on_commit : _GEN_6467
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6666 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_unique : _GEN_6468; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6667 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_sys_pc2epc : _GEN_6469; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6668 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_uses_stq : _GEN_6470; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6669 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_uses_ldq : _GEN_6471; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6670 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_amo : _GEN_6472; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6671 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_fencei : _GEN_6473; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6672 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_fence : _GEN_6474; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6673 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_mem_signed : _GEN_6475; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6674 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_mem_size : _GEN_6476; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6675 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_mem_cmd : _GEN_6477; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6676 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_bypassable : _GEN_6478; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_6677 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_exc_cause : _GEN_6479
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6678 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_exception : _GEN_6480; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6679 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_stale_pdst : _GEN_6481
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6680 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ppred_busy : _GEN_6482; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6681 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_prs3_busy : _GEN_6483; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6682 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_prs2_busy : _GEN_6484; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6683 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_prs1_busy : _GEN_6485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6684 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ppred : _GEN_6486; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6685 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_prs3 : _GEN_6487; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6686 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_prs2 : _GEN_6488; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6687 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_prs1 : _GEN_6489; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6688 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_pdst : _GEN_6490; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6689 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_rxq_idx : _GEN_6491; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6690 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_stq_idx : _GEN_6492; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6691 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ldq_idx : _GEN_6493; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6692 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_rob_idx : _GEN_6494; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6693 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_csr_addr : _GEN_6495; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_6694 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_imm_packed :
    _GEN_6496; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6695 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_taken : _GEN_6497; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6696 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_pc_lob : _GEN_6498; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6697 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_edge_inst : _GEN_6499; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6698 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ftq_idx : _GEN_6500; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6699 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_br_tag : _GEN_6501; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6700 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_br_mask : _GEN_6502; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6701 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_sfb : _GEN_6503; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6702 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_jal : _GEN_6504; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6703 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_jalr : _GEN_6505; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6704 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_br : _GEN_6506; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6705 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_iw_p2_poisoned : _GEN_6507; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6706 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_iw_p1_poisoned : _GEN_6508; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6707 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_iw_state : _GEN_6509; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6708 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_op3_sel :
    _GEN_6510; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6709 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_is_std : _GEN_6511; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6710 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_is_sta : _GEN_6512; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6711 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_is_load : _GEN_6513; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6712 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_csr_cmd :
    _GEN_6514; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6713 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_fcn_dw : _GEN_6515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6714 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_op_fcn :
    _GEN_6516; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6715 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_imm_sel :
    _GEN_6517; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6716 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_op2_sel :
    _GEN_6518; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6717 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_op1_sel :
    _GEN_6519; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6718 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_ctrl_br_type :
    _GEN_6520; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6719 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_fu_code : _GEN_6521; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6720 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_iq_type : _GEN_6522; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_6721 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_debug_pc : _GEN_6523; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6722 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_rvc : _GEN_6524; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6723 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_debug_inst :
    _GEN_6525; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6724 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_inst : _GEN_6526; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6725 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_uopc : _GEN_6527; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6726 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_address_num :
    _GEN_6528; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6727 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_rob_inst_idx :
    _GEN_6529; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6728 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_self_index : _GEN_6530
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6729 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_split_num : _GEN_6531; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6730 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_op2_sel : _GEN_6532; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6731 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_op1_sel : _GEN_6533; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6732 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_stale_pflag :
    _GEN_6534; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6733 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_pflag_busy : _GEN_6535; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6734 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_pwflag : _GEN_6536; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6735 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_prflag : _GEN_6537; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6736 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_wflag : _GEN_6538; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6737 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_rflag : _GEN_6539; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6738 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_lrs3_rtype : _GEN_6540
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6739 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_shift : _GEN_6541; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6740 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_is_unicore : _GEN_6542; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6741 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_switch_off : _GEN_6543; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6742 = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 ? issue_slots_13_uop_switch : _GEN_6544; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_debug_tsrc = slots_14_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6745 = _T_845 ? issue_slots_14_uop_debug_tsrc : _GEN_6547; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_debug_fsrc = slots_14_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6746 = _T_845 ? issue_slots_14_uop_debug_fsrc : _GEN_6548; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_bp_xcpt_if = slots_14_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6747 = _T_845 ? issue_slots_14_uop_bp_xcpt_if : _GEN_6549; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_bp_debug_if = slots_14_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6748 = _T_845 ? issue_slots_14_uop_bp_debug_if : _GEN_6550; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_xcpt_ma_if = slots_14_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6749 = _T_845 ? issue_slots_14_uop_xcpt_ma_if : _GEN_6551; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_xcpt_ae_if = slots_14_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6750 = _T_845 ? issue_slots_14_uop_xcpt_ae_if : _GEN_6552; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_xcpt_pf_if = slots_14_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6751 = _T_845 ? issue_slots_14_uop_xcpt_pf_if : _GEN_6553; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_fp_single = slots_14_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6752 = _T_845 ? issue_slots_14_uop_fp_single : _GEN_6554; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_fp_val = slots_14_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6753 = _T_845 ? issue_slots_14_uop_fp_val : _GEN_6555; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_frs3_en = slots_14_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6754 = _T_845 ? issue_slots_14_uop_frs3_en : _GEN_6556; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_lrs2_rtype = slots_14_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6755 = _T_845 ? issue_slots_14_uop_lrs2_rtype : _GEN_6557; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_lrs1_rtype = slots_14_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6756 = _T_845 ? issue_slots_14_uop_lrs1_rtype : _GEN_6558; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_dst_rtype = slots_14_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6757 = _T_845 ? issue_slots_14_uop_dst_rtype : _GEN_6559; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ldst_val = slots_14_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6758 = _T_845 ? issue_slots_14_uop_ldst_val : _GEN_6560; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_lrs3 = slots_14_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6759 = _T_845 ? issue_slots_14_uop_lrs3 : _GEN_6561; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_lrs2 = slots_14_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6760 = _T_845 ? issue_slots_14_uop_lrs2 : _GEN_6562; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_lrs1 = slots_14_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6761 = _T_845 ? issue_slots_14_uop_lrs1 : _GEN_6563; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_ldst = slots_14_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6762 = _T_845 ? issue_slots_14_uop_ldst : _GEN_6564; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ldst_is_rs1 = slots_14_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6763 = _T_845 ? issue_slots_14_uop_ldst_is_rs1 : _GEN_6565; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_flush_on_commit = slots_14_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6764 = _T_845 ? issue_slots_14_uop_flush_on_commit : _GEN_6566; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_unique = slots_14_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6765 = _T_845 ? issue_slots_14_uop_is_unique : _GEN_6567; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_sys_pc2epc = slots_14_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6766 = _T_845 ? issue_slots_14_uop_is_sys_pc2epc : _GEN_6568; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_uses_stq = slots_14_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6767 = _T_845 ? issue_slots_14_uop_uses_stq : _GEN_6569; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_uses_ldq = slots_14_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6768 = _T_845 ? issue_slots_14_uop_uses_ldq : _GEN_6570; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_amo = slots_14_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6769 = _T_845 ? issue_slots_14_uop_is_amo : _GEN_6571; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_fencei = slots_14_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6770 = _T_845 ? issue_slots_14_uop_is_fencei : _GEN_6572; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_fence = slots_14_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6771 = _T_845 ? issue_slots_14_uop_is_fence : _GEN_6573; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_mem_signed = slots_14_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6772 = _T_845 ? issue_slots_14_uop_mem_signed : _GEN_6574; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_mem_size = slots_14_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6773 = _T_845 ? issue_slots_14_uop_mem_size : _GEN_6575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_mem_cmd = slots_14_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6774 = _T_845 ? issue_slots_14_uop_mem_cmd : _GEN_6576; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_bypassable = slots_14_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6775 = _T_845 ? issue_slots_14_uop_bypassable : _GEN_6577; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_14_uop_exc_cause = slots_14_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_6776 = _T_845 ? issue_slots_14_uop_exc_cause : _GEN_6578; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_exception = slots_14_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6777 = _T_845 ? issue_slots_14_uop_exception : _GEN_6579; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_stale_pdst = slots_14_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6778 = _T_845 ? issue_slots_14_uop_stale_pdst : _GEN_6580; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ppred_busy = slots_14_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6779 = _T_845 ? issue_slots_14_uop_ppred_busy : _GEN_6581; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_prs3_busy = slots_14_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6780 = _T_845 ? issue_slots_14_uop_prs3_busy : _GEN_6582; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_prs2_busy = slots_14_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6781 = _T_845 ? issue_slots_14_uop_prs2_busy : _GEN_6583; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_prs1_busy = slots_14_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6782 = _T_845 ? issue_slots_14_uop_prs1_busy : _GEN_6584; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_ppred = slots_14_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6783 = _T_845 ? issue_slots_14_uop_ppred : _GEN_6585; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_prs3 = slots_14_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6784 = _T_845 ? issue_slots_14_uop_prs3 : _GEN_6586; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_prs2 = slots_14_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6785 = _T_845 ? issue_slots_14_uop_prs2 : _GEN_6587; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_prs1 = slots_14_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6786 = _T_845 ? issue_slots_14_uop_prs1 : _GEN_6588; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_pdst = slots_14_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6787 = _T_845 ? issue_slots_14_uop_pdst : _GEN_6589; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_rxq_idx = slots_14_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6788 = _T_845 ? issue_slots_14_uop_rxq_idx : _GEN_6590; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_stq_idx = slots_14_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6789 = _T_845 ? issue_slots_14_uop_stq_idx : _GEN_6591; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_ldq_idx = slots_14_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6790 = _T_845 ? issue_slots_14_uop_ldq_idx : _GEN_6592; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_rob_idx = slots_14_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6791 = _T_845 ? issue_slots_14_uop_rob_idx : _GEN_6593; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_14_uop_csr_addr = slots_14_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6792 = _T_845 ? issue_slots_14_uop_csr_addr : _GEN_6594; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_14_uop_imm_packed = slots_14_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_6793 = _T_845 ? issue_slots_14_uop_imm_packed : _GEN_6595; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_taken = slots_14_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6794 = _T_845 ? issue_slots_14_uop_taken : _GEN_6596; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_pc_lob = slots_14_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6795 = _T_845 ? issue_slots_14_uop_pc_lob : _GEN_6597; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_edge_inst = slots_14_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6796 = _T_845 ? issue_slots_14_uop_edge_inst : _GEN_6598; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_ftq_idx = slots_14_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6797 = _T_845 ? issue_slots_14_uop_ftq_idx : _GEN_6599; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_br_tag = slots_14_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6798 = _T_845 ? issue_slots_14_uop_br_tag : _GEN_6600; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_14_uop_br_mask = slots_14_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6799 = _T_845 ? issue_slots_14_uop_br_mask : _GEN_6601; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_sfb = slots_14_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6800 = _T_845 ? issue_slots_14_uop_is_sfb : _GEN_6602; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_jal = slots_14_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6801 = _T_845 ? issue_slots_14_uop_is_jal : _GEN_6603; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_jalr = slots_14_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6802 = _T_845 ? issue_slots_14_uop_is_jalr : _GEN_6604; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_br = slots_14_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6803 = _T_845 ? issue_slots_14_uop_is_br : _GEN_6605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_iw_p2_poisoned = slots_14_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6804 = _T_845 ? issue_slots_14_uop_iw_p2_poisoned : _GEN_6606; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_iw_p1_poisoned = slots_14_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6805 = _T_845 ? issue_slots_14_uop_iw_p1_poisoned : _GEN_6607; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_iw_state = slots_14_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6806 = _T_845 ? issue_slots_14_uop_iw_state : _GEN_6608; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_ctrl_op3_sel = slots_14_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6807 = _T_845 ? issue_slots_14_uop_ctrl_op3_sel : _GEN_6609; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_is_std = slots_14_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6808 = _T_845 ? issue_slots_14_uop_ctrl_is_std : _GEN_6610; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_is_sta = slots_14_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6809 = _T_845 ? issue_slots_14_uop_ctrl_is_sta : _GEN_6611; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_is_load = slots_14_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6810 = _T_845 ? issue_slots_14_uop_ctrl_is_load : _GEN_6612; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_ctrl_csr_cmd = slots_14_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6811 = _T_845 ? issue_slots_14_uop_ctrl_csr_cmd : _GEN_6613; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_fcn_dw = slots_14_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6812 = _T_845 ? issue_slots_14_uop_ctrl_fcn_dw : _GEN_6614; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_ctrl_op_fcn = slots_14_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6813 = _T_845 ? issue_slots_14_uop_ctrl_op_fcn : _GEN_6615; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_ctrl_imm_sel = slots_14_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6814 = _T_845 ? issue_slots_14_uop_ctrl_imm_sel : _GEN_6616; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_ctrl_op2_sel = slots_14_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6815 = _T_845 ? issue_slots_14_uop_ctrl_op2_sel : _GEN_6617; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_ctrl_op1_sel = slots_14_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6816 = _T_845 ? issue_slots_14_uop_ctrl_op1_sel : _GEN_6618; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_ctrl_br_type = slots_14_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6817 = _T_845 ? issue_slots_14_uop_ctrl_br_type : _GEN_6619; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6818 = _T_845 ? issue_slots_14_uop_fu_code : _GEN_6620; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_iq_type = slots_14_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6819 = _T_845 ? issue_slots_14_uop_iq_type : _GEN_6621; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_14_uop_debug_pc = slots_14_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_6820 = _T_845 ? issue_slots_14_uop_debug_pc : _GEN_6622; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_rvc = slots_14_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6821 = _T_845 ? issue_slots_14_uop_is_rvc : _GEN_6623; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_14_uop_debug_inst = slots_14_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6822 = _T_845 ? issue_slots_14_uop_debug_inst : _GEN_6624; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_14_uop_inst = slots_14_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_6823 = _T_845 ? issue_slots_14_uop_inst : _GEN_6625; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_uopc = slots_14_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6824 = _T_845 ? issue_slots_14_uop_uopc : _GEN_6626; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_address_num = slots_14_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6825 = _T_845 ? issue_slots_14_uop_address_num : _GEN_6627; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_rob_inst_idx = slots_14_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6826 = _T_845 ? issue_slots_14_uop_rob_inst_idx : _GEN_6628; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_self_index = slots_14_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6827 = _T_845 ? issue_slots_14_uop_self_index : _GEN_6629; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_split_num = slots_14_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6828 = _T_845 ? issue_slots_14_uop_split_num : _GEN_6630; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_op2_sel = slots_14_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6829 = _T_845 ? issue_slots_14_uop_op2_sel : _GEN_6631; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_op1_sel = slots_14_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6830 = _T_845 ? issue_slots_14_uop_op1_sel : _GEN_6632; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_stale_pflag = slots_14_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6831 = _T_845 ? issue_slots_14_uop_stale_pflag : _GEN_6633; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_pflag_busy = slots_14_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6832 = _T_845 ? issue_slots_14_uop_pflag_busy : _GEN_6634; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_pwflag = slots_14_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6833 = _T_845 ? issue_slots_14_uop_pwflag : _GEN_6635; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_prflag = slots_14_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6834 = _T_845 ? issue_slots_14_uop_prflag : _GEN_6636; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_wflag = slots_14_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6835 = _T_845 ? issue_slots_14_uop_wflag : _GEN_6637; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_rflag = slots_14_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6836 = _T_845 ? issue_slots_14_uop_rflag : _GEN_6638; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_lrs3_rtype = slots_14_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6837 = _T_845 ? issue_slots_14_uop_lrs3_rtype : _GEN_6639; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_shift = slots_14_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_6838 = _T_845 ? issue_slots_14_uop_shift : _GEN_6640; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_unicore = slots_14_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6839 = _T_845 ? issue_slots_14_uop_is_unicore : _GEN_6641; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_switch_off = slots_14_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6840 = _T_845 ? issue_slots_14_uop_switch_off : _GEN_6642; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_switch = slots_14_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6841 = _T_845 ? issue_slots_14_uop_switch : _GEN_6643; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6843 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 | (issue_slots_13_request & ~_T_815 & _T_818 & ~
    _T_797 | (_T_796 & ~_T_767 | (issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 | (issue_slots_10_request & ~
    _T_725 & _T_728 & ~_T_707 | _GEN_5853)))); // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 124:26]
  wire [1:0] _GEN_6844 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_debug_tsrc : _GEN_6646
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6845 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_debug_fsrc : _GEN_6647
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6846 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_bp_xcpt_if : _GEN_6648; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6847 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_bp_debug_if : _GEN_6649; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6848 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_xcpt_ma_if : _GEN_6650; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6849 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_xcpt_ae_if : _GEN_6651; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6850 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_xcpt_pf_if : _GEN_6652; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6851 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_fp_single : _GEN_6653; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6852 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_fp_val : _GEN_6654; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6853 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_frs3_en : _GEN_6655; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6854 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_lrs2_rtype : _GEN_6656
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6855 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_lrs1_rtype : _GEN_6657
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6856 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_dst_rtype : _GEN_6658; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6857 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ldst_val : _GEN_6659; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6858 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_lrs3 : _GEN_6660; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6859 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_lrs2 : _GEN_6661; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6860 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_lrs1 : _GEN_6662; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6861 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ldst : _GEN_6663; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6862 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ldst_is_rs1 : _GEN_6664; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6863 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_flush_on_commit : _GEN_6665
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6864 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_unique : _GEN_6666; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6865 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_sys_pc2epc : _GEN_6667; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6866 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_uses_stq : _GEN_6668; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6867 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_uses_ldq : _GEN_6669; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6868 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_amo : _GEN_6670; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6869 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_fencei : _GEN_6671; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6870 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_fence : _GEN_6672; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6871 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_mem_signed : _GEN_6673; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6872 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_mem_size : _GEN_6674; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6873 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_mem_cmd : _GEN_6675; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6874 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_bypassable : _GEN_6676; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_6875 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_exc_cause : _GEN_6677
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6876 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_exception : _GEN_6678; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6877 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_stale_pdst : _GEN_6679
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6878 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ppred_busy : _GEN_6680; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6879 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_prs3_busy : _GEN_6681; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6880 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_prs2_busy : _GEN_6682; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6881 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_prs1_busy : _GEN_6683; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6882 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ppred : _GEN_6684; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6883 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_prs3 : _GEN_6685; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6884 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_prs2 : _GEN_6686; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6885 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_prs1 : _GEN_6687; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6886 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_pdst : _GEN_6688; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6887 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_rxq_idx : _GEN_6689; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6888 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_stq_idx : _GEN_6690; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6889 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ldq_idx : _GEN_6691; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6890 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_rob_idx : _GEN_6692; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6891 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_csr_addr : _GEN_6693; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_6892 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_imm_packed :
    _GEN_6694; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6893 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_taken : _GEN_6695; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6894 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_pc_lob : _GEN_6696; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6895 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_edge_inst : _GEN_6697; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_6896 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ftq_idx : _GEN_6698; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6897 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_br_tag : _GEN_6699; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_6898 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_br_mask : _GEN_6700; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6899 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_sfb : _GEN_6701; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6900 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_jal : _GEN_6702; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6901 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_jalr : _GEN_6703; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6902 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_br : _GEN_6704; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6903 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_iw_p2_poisoned : _GEN_6705; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6904 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_iw_p1_poisoned : _GEN_6706; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6905 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_iw_state : _GEN_6707; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6906 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_op3_sel :
    _GEN_6708; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6907 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_is_std : _GEN_6709; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6908 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_is_sta : _GEN_6710; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6909 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_is_load : _GEN_6711; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6910 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_csr_cmd :
    _GEN_6712; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6911 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_fcn_dw : _GEN_6713; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6912 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_op_fcn :
    _GEN_6714; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6913 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_imm_sel :
    _GEN_6715; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6914 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_op2_sel :
    _GEN_6716; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6915 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_op1_sel :
    _GEN_6717; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6916 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_ctrl_br_type :
    _GEN_6718; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_6917 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_fu_code : _GEN_6719; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6918 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_iq_type : _GEN_6720; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_6919 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_debug_pc : _GEN_6721; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6920 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_rvc : _GEN_6722; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6921 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_debug_inst :
    _GEN_6723; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_6922 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_inst : _GEN_6724; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_6923 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_uopc : _GEN_6725; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6924 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_address_num :
    _GEN_6726; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6925 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_rob_inst_idx :
    _GEN_6727; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6926 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_self_index : _GEN_6728
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_6927 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_split_num : _GEN_6729; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6928 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_op2_sel : _GEN_6730; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6929 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_op1_sel : _GEN_6731; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6930 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_stale_pflag :
    _GEN_6732; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6931 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_pflag_busy : _GEN_6733; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6932 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_pwflag : _GEN_6734; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_6933 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_prflag : _GEN_6735; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6934 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_wflag : _GEN_6736; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6935 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_rflag : _GEN_6737; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_6936 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_lrs3_rtype : _GEN_6738
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_6937 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_shift : _GEN_6739; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6938 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_is_unicore : _GEN_6740; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6939 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_switch_off : _GEN_6741; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_6940 = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 ? issue_slots_14_uop_switch : _GEN_6742; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_debug_tsrc = slots_15_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6943 = _T_875 ? issue_slots_15_uop_debug_tsrc : _GEN_6745; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_debug_fsrc = slots_15_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6944 = _T_875 ? issue_slots_15_uop_debug_fsrc : _GEN_6746; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_bp_xcpt_if = slots_15_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6945 = _T_875 ? issue_slots_15_uop_bp_xcpt_if : _GEN_6747; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_bp_debug_if = slots_15_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6946 = _T_875 ? issue_slots_15_uop_bp_debug_if : _GEN_6748; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_xcpt_ma_if = slots_15_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6947 = _T_875 ? issue_slots_15_uop_xcpt_ma_if : _GEN_6749; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_xcpt_ae_if = slots_15_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6948 = _T_875 ? issue_slots_15_uop_xcpt_ae_if : _GEN_6750; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_xcpt_pf_if = slots_15_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6949 = _T_875 ? issue_slots_15_uop_xcpt_pf_if : _GEN_6751; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_fp_single = slots_15_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6950 = _T_875 ? issue_slots_15_uop_fp_single : _GEN_6752; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_fp_val = slots_15_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6951 = _T_875 ? issue_slots_15_uop_fp_val : _GEN_6753; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_frs3_en = slots_15_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6952 = _T_875 ? issue_slots_15_uop_frs3_en : _GEN_6754; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_lrs2_rtype = slots_15_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6953 = _T_875 ? issue_slots_15_uop_lrs2_rtype : _GEN_6755; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_lrs1_rtype = slots_15_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6954 = _T_875 ? issue_slots_15_uop_lrs1_rtype : _GEN_6756; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_dst_rtype = slots_15_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6955 = _T_875 ? issue_slots_15_uop_dst_rtype : _GEN_6757; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_ldst_val = slots_15_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6956 = _T_875 ? issue_slots_15_uop_ldst_val : _GEN_6758; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_lrs3 = slots_15_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6957 = _T_875 ? issue_slots_15_uop_lrs3 : _GEN_6759; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_lrs2 = slots_15_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6958 = _T_875 ? issue_slots_15_uop_lrs2 : _GEN_6760; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_lrs1 = slots_15_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6959 = _T_875 ? issue_slots_15_uop_lrs1 : _GEN_6761; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_ldst = slots_15_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6960 = _T_875 ? issue_slots_15_uop_ldst : _GEN_6762; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_ldst_is_rs1 = slots_15_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6961 = _T_875 ? issue_slots_15_uop_ldst_is_rs1 : _GEN_6763; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_flush_on_commit = slots_15_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6962 = _T_875 ? issue_slots_15_uop_flush_on_commit : _GEN_6764; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_unique = slots_15_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6963 = _T_875 ? issue_slots_15_uop_is_unique : _GEN_6765; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_sys_pc2epc = slots_15_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6964 = _T_875 ? issue_slots_15_uop_is_sys_pc2epc : _GEN_6766; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_uses_stq = slots_15_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6965 = _T_875 ? issue_slots_15_uop_uses_stq : _GEN_6767; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_uses_ldq = slots_15_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6966 = _T_875 ? issue_slots_15_uop_uses_ldq : _GEN_6768; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_amo = slots_15_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6967 = _T_875 ? issue_slots_15_uop_is_amo : _GEN_6769; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_fencei = slots_15_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6968 = _T_875 ? issue_slots_15_uop_is_fencei : _GEN_6770; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_fence = slots_15_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6969 = _T_875 ? issue_slots_15_uop_is_fence : _GEN_6771; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_mem_signed = slots_15_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6970 = _T_875 ? issue_slots_15_uop_mem_signed : _GEN_6772; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_mem_size = slots_15_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6971 = _T_875 ? issue_slots_15_uop_mem_size : _GEN_6773; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_15_uop_mem_cmd = slots_15_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6972 = _T_875 ? issue_slots_15_uop_mem_cmd : _GEN_6774; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_bypassable = slots_15_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6973 = _T_875 ? issue_slots_15_uop_bypassable : _GEN_6775; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_15_uop_exc_cause = slots_15_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_6974 = _T_875 ? issue_slots_15_uop_exc_cause : _GEN_6776; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_exception = slots_15_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6975 = _T_875 ? issue_slots_15_uop_exception : _GEN_6777; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_15_uop_stale_pdst = slots_15_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6976 = _T_875 ? issue_slots_15_uop_stale_pdst : _GEN_6778; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_ppred_busy = slots_15_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6977 = _T_875 ? issue_slots_15_uop_ppred_busy : _GEN_6779; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_prs3_busy = slots_15_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6978 = _T_875 ? issue_slots_15_uop_prs3_busy : _GEN_6780; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_prs2_busy = slots_15_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6979 = _T_875 ? issue_slots_15_uop_prs2_busy : _GEN_6781; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_prs1_busy = slots_15_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6980 = _T_875 ? issue_slots_15_uop_prs1_busy : _GEN_6782; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_15_uop_ppred = slots_15_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6981 = _T_875 ? issue_slots_15_uop_ppred : _GEN_6783; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_15_uop_prs3 = slots_15_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6982 = _T_875 ? issue_slots_15_uop_prs3 : _GEN_6784; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_15_uop_prs2 = slots_15_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6983 = _T_875 ? issue_slots_15_uop_prs2 : _GEN_6785; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_15_uop_prs1 = slots_15_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6984 = _T_875 ? issue_slots_15_uop_prs1 : _GEN_6786; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_15_uop_pdst = slots_15_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_6985 = _T_875 ? issue_slots_15_uop_pdst : _GEN_6787; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_rxq_idx = slots_15_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_6986 = _T_875 ? issue_slots_15_uop_rxq_idx : _GEN_6788; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_15_uop_stq_idx = slots_15_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6987 = _T_875 ? issue_slots_15_uop_stq_idx : _GEN_6789; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_15_uop_ldq_idx = slots_15_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6988 = _T_875 ? issue_slots_15_uop_ldq_idx : _GEN_6790; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_rob_idx = slots_15_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6989 = _T_875 ? issue_slots_15_uop_rob_idx : _GEN_6791; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_15_uop_csr_addr = slots_15_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6990 = _T_875 ? issue_slots_15_uop_csr_addr : _GEN_6792; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_15_uop_imm_packed = slots_15_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_6991 = _T_875 ? issue_slots_15_uop_imm_packed : _GEN_6793; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_taken = slots_15_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6992 = _T_875 ? issue_slots_15_uop_taken : _GEN_6794; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_pc_lob = slots_15_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_6993 = _T_875 ? issue_slots_15_uop_pc_lob : _GEN_6795; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_edge_inst = slots_15_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6994 = _T_875 ? issue_slots_15_uop_edge_inst : _GEN_6796; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_15_uop_ftq_idx = slots_15_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_6995 = _T_875 ? issue_slots_15_uop_ftq_idx : _GEN_6797; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_br_tag = slots_15_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_6996 = _T_875 ? issue_slots_15_uop_br_tag : _GEN_6798; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_15_uop_br_mask = slots_15_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_6997 = _T_875 ? issue_slots_15_uop_br_mask : _GEN_6799; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_sfb = slots_15_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6998 = _T_875 ? issue_slots_15_uop_is_sfb : _GEN_6800; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_jal = slots_15_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_6999 = _T_875 ? issue_slots_15_uop_is_jal : _GEN_6801; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_jalr = slots_15_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7000 = _T_875 ? issue_slots_15_uop_is_jalr : _GEN_6802; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_br = slots_15_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7001 = _T_875 ? issue_slots_15_uop_is_br : _GEN_6803; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_iw_p2_poisoned = slots_15_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7002 = _T_875 ? issue_slots_15_uop_iw_p2_poisoned : _GEN_6804; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_iw_p1_poisoned = slots_15_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7003 = _T_875 ? issue_slots_15_uop_iw_p1_poisoned : _GEN_6805; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_iw_state = slots_15_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7004 = _T_875 ? issue_slots_15_uop_iw_state : _GEN_6806; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_ctrl_op3_sel = slots_15_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7005 = _T_875 ? issue_slots_15_uop_ctrl_op3_sel : _GEN_6807; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_ctrl_is_std = slots_15_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7006 = _T_875 ? issue_slots_15_uop_ctrl_is_std : _GEN_6808; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_ctrl_is_sta = slots_15_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7007 = _T_875 ? issue_slots_15_uop_ctrl_is_sta : _GEN_6809; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_ctrl_is_load = slots_15_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7008 = _T_875 ? issue_slots_15_uop_ctrl_is_load : _GEN_6810; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_15_uop_ctrl_csr_cmd = slots_15_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7009 = _T_875 ? issue_slots_15_uop_ctrl_csr_cmd : _GEN_6811; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_ctrl_fcn_dw = slots_15_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7010 = _T_875 ? issue_slots_15_uop_ctrl_fcn_dw : _GEN_6812; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_ctrl_op_fcn = slots_15_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7011 = _T_875 ? issue_slots_15_uop_ctrl_op_fcn : _GEN_6813; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_15_uop_ctrl_imm_sel = slots_15_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7012 = _T_875 ? issue_slots_15_uop_ctrl_imm_sel : _GEN_6814; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_15_uop_ctrl_op2_sel = slots_15_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7013 = _T_875 ? issue_slots_15_uop_ctrl_op2_sel : _GEN_6815; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_ctrl_op1_sel = slots_15_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7014 = _T_875 ? issue_slots_15_uop_ctrl_op1_sel : _GEN_6816; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_ctrl_br_type = slots_15_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7015 = _T_875 ? issue_slots_15_uop_ctrl_br_type : _GEN_6817; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7016 = _T_875 ? issue_slots_15_uop_fu_code : _GEN_6818; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_15_uop_iq_type = slots_15_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7017 = _T_875 ? issue_slots_15_uop_iq_type : _GEN_6819; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_15_uop_debug_pc = slots_15_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_7018 = _T_875 ? issue_slots_15_uop_debug_pc : _GEN_6820; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_rvc = slots_15_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7019 = _T_875 ? issue_slots_15_uop_is_rvc : _GEN_6821; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_15_uop_debug_inst = slots_15_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7020 = _T_875 ? issue_slots_15_uop_debug_inst : _GEN_6822; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_15_uop_inst = slots_15_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7021 = _T_875 ? issue_slots_15_uop_inst : _GEN_6823; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_15_uop_uopc = slots_15_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7022 = _T_875 ? issue_slots_15_uop_uopc : _GEN_6824; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_address_num = slots_15_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7023 = _T_875 ? issue_slots_15_uop_address_num : _GEN_6825; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_rob_inst_idx = slots_15_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7024 = _T_875 ? issue_slots_15_uop_rob_inst_idx : _GEN_6826; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_self_index = slots_15_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7025 = _T_875 ? issue_slots_15_uop_self_index : _GEN_6827; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_15_uop_split_num = slots_15_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7026 = _T_875 ? issue_slots_15_uop_split_num : _GEN_6828; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_op2_sel = slots_15_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7027 = _T_875 ? issue_slots_15_uop_op2_sel : _GEN_6829; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_op1_sel = slots_15_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7028 = _T_875 ? issue_slots_15_uop_op1_sel : _GEN_6830; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_stale_pflag = slots_15_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7029 = _T_875 ? issue_slots_15_uop_stale_pflag : _GEN_6831; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_pflag_busy = slots_15_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7030 = _T_875 ? issue_slots_15_uop_pflag_busy : _GEN_6832; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_pwflag = slots_15_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7031 = _T_875 ? issue_slots_15_uop_pwflag : _GEN_6833; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_15_uop_prflag = slots_15_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7032 = _T_875 ? issue_slots_15_uop_prflag : _GEN_6834; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_wflag = slots_15_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7033 = _T_875 ? issue_slots_15_uop_wflag : _GEN_6835; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_rflag = slots_15_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7034 = _T_875 ? issue_slots_15_uop_rflag : _GEN_6836; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_lrs3_rtype = slots_15_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7035 = _T_875 ? issue_slots_15_uop_lrs3_rtype : _GEN_6837; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_15_uop_shift = slots_15_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7036 = _T_875 ? issue_slots_15_uop_shift : _GEN_6838; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_is_unicore = slots_15_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7037 = _T_875 ? issue_slots_15_uop_is_unicore : _GEN_6839; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_switch_off = slots_15_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7038 = _T_875 ? issue_slots_15_uop_switch_off : _GEN_6840; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_15_uop_switch = slots_15_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7039 = _T_875 ? issue_slots_15_uop_switch : _GEN_6841; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7042 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_debug_tsrc : _GEN_6844
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7043 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_debug_fsrc : _GEN_6845
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7044 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_bp_xcpt_if : _GEN_6846; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7045 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_bp_debug_if : _GEN_6847; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7046 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_xcpt_ma_if : _GEN_6848; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7047 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_xcpt_ae_if : _GEN_6849; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7048 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_xcpt_pf_if : _GEN_6850; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7049 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_fp_single : _GEN_6851; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7050 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_fp_val : _GEN_6852; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7051 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_frs3_en : _GEN_6853; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7052 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_lrs2_rtype : _GEN_6854
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7053 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_lrs1_rtype : _GEN_6855
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7054 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_dst_rtype : _GEN_6856; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7055 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ldst_val : _GEN_6857; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7056 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_lrs3 : _GEN_6858; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7057 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_lrs2 : _GEN_6859; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7058 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_lrs1 : _GEN_6860; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7059 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ldst : _GEN_6861; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7060 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ldst_is_rs1 : _GEN_6862; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7061 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_flush_on_commit : _GEN_6863
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7062 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_unique : _GEN_6864; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7063 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_sys_pc2epc : _GEN_6865; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7064 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_uses_stq : _GEN_6866; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7065 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_uses_ldq : _GEN_6867; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7066 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_amo : _GEN_6868; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7067 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_fencei : _GEN_6869; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7068 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_fence : _GEN_6870; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7069 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_mem_signed : _GEN_6871; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7070 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_mem_size : _GEN_6872; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7071 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_mem_cmd : _GEN_6873; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7072 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_bypassable : _GEN_6874; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_7073 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_exc_cause : _GEN_6875
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7074 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_exception : _GEN_6876; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7075 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_stale_pdst : _GEN_6877
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7076 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ppred_busy : _GEN_6878; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7077 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_prs3_busy : _GEN_6879; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7078 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_prs2_busy : _GEN_6880; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7079 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_prs1_busy : _GEN_6881; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7080 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ppred : _GEN_6882; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7081 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_prs3 : _GEN_6883; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7082 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_prs2 : _GEN_6884; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7083 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_prs1 : _GEN_6885; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7084 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_pdst : _GEN_6886; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7085 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_rxq_idx : _GEN_6887; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7086 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_stq_idx : _GEN_6888; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7087 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ldq_idx : _GEN_6889; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7088 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_rob_idx : _GEN_6890; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7089 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_csr_addr : _GEN_6891; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_7090 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_imm_packed :
    _GEN_6892; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7091 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_taken : _GEN_6893; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7092 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_pc_lob : _GEN_6894; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7093 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_edge_inst : _GEN_6895; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7094 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ftq_idx : _GEN_6896; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7095 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_br_tag : _GEN_6897; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7096 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_br_mask : _GEN_6898; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7097 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_sfb : _GEN_6899; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7098 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_jal : _GEN_6900; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7099 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_jalr : _GEN_6901; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7100 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_br : _GEN_6902; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7101 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_iw_p2_poisoned : _GEN_6903; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7102 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_iw_p1_poisoned : _GEN_6904; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7103 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_iw_state : _GEN_6905; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7104 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_op3_sel :
    _GEN_6906; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7105 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_is_std : _GEN_6907; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7106 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_is_sta : _GEN_6908; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7107 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_is_load : _GEN_6909; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7108 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_csr_cmd :
    _GEN_6910; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7109 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_fcn_dw : _GEN_6911; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7110 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_op_fcn :
    _GEN_6912; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7111 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_imm_sel :
    _GEN_6913; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7112 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_op2_sel :
    _GEN_6914; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7113 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_op1_sel :
    _GEN_6915; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7114 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_ctrl_br_type :
    _GEN_6916; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7115 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_fu_code : _GEN_6917; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7116 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_iq_type : _GEN_6918; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_7117 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_debug_pc : _GEN_6919; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7118 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_rvc : _GEN_6920; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7119 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_debug_inst :
    _GEN_6921; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7120 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_inst : _GEN_6922; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7121 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_uopc : _GEN_6923; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7122 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_address_num :
    _GEN_6924; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7123 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_rob_inst_idx :
    _GEN_6925; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7124 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_self_index : _GEN_6926
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7125 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_split_num : _GEN_6927; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7126 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_op2_sel : _GEN_6928; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7127 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_op1_sel : _GEN_6929; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7128 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_stale_pflag :
    _GEN_6930; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7129 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_pflag_busy : _GEN_6931; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7130 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_pwflag : _GEN_6932; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7131 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_prflag : _GEN_6933; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7132 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_wflag : _GEN_6934; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7133 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_rflag : _GEN_6935; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7134 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_lrs3_rtype : _GEN_6936
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7135 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_shift : _GEN_6937; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7136 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_is_unicore : _GEN_6938; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7137 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_switch_off : _GEN_6939; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7138 = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 ? issue_slots_15_uop_switch : _GEN_6940; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_debug_tsrc = slots_16_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7141 = _T_905 ? issue_slots_16_uop_debug_tsrc : _GEN_6943; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_debug_fsrc = slots_16_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7142 = _T_905 ? issue_slots_16_uop_debug_fsrc : _GEN_6944; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_bp_xcpt_if = slots_16_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7143 = _T_905 ? issue_slots_16_uop_bp_xcpt_if : _GEN_6945; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_bp_debug_if = slots_16_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7144 = _T_905 ? issue_slots_16_uop_bp_debug_if : _GEN_6946; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_xcpt_ma_if = slots_16_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7145 = _T_905 ? issue_slots_16_uop_xcpt_ma_if : _GEN_6947; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_xcpt_ae_if = slots_16_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7146 = _T_905 ? issue_slots_16_uop_xcpt_ae_if : _GEN_6948; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_xcpt_pf_if = slots_16_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7147 = _T_905 ? issue_slots_16_uop_xcpt_pf_if : _GEN_6949; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_fp_single = slots_16_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7148 = _T_905 ? issue_slots_16_uop_fp_single : _GEN_6950; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_fp_val = slots_16_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7149 = _T_905 ? issue_slots_16_uop_fp_val : _GEN_6951; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_frs3_en = slots_16_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7150 = _T_905 ? issue_slots_16_uop_frs3_en : _GEN_6952; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_lrs2_rtype = slots_16_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7151 = _T_905 ? issue_slots_16_uop_lrs2_rtype : _GEN_6953; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_lrs1_rtype = slots_16_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7152 = _T_905 ? issue_slots_16_uop_lrs1_rtype : _GEN_6954; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_dst_rtype = slots_16_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7153 = _T_905 ? issue_slots_16_uop_dst_rtype : _GEN_6955; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_ldst_val = slots_16_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7154 = _T_905 ? issue_slots_16_uop_ldst_val : _GEN_6956; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_lrs3 = slots_16_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7155 = _T_905 ? issue_slots_16_uop_lrs3 : _GEN_6957; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_lrs2 = slots_16_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7156 = _T_905 ? issue_slots_16_uop_lrs2 : _GEN_6958; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_lrs1 = slots_16_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7157 = _T_905 ? issue_slots_16_uop_lrs1 : _GEN_6959; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_ldst = slots_16_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7158 = _T_905 ? issue_slots_16_uop_ldst : _GEN_6960; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_ldst_is_rs1 = slots_16_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7159 = _T_905 ? issue_slots_16_uop_ldst_is_rs1 : _GEN_6961; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_flush_on_commit = slots_16_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7160 = _T_905 ? issue_slots_16_uop_flush_on_commit : _GEN_6962; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_unique = slots_16_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7161 = _T_905 ? issue_slots_16_uop_is_unique : _GEN_6963; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_sys_pc2epc = slots_16_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7162 = _T_905 ? issue_slots_16_uop_is_sys_pc2epc : _GEN_6964; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_uses_stq = slots_16_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7163 = _T_905 ? issue_slots_16_uop_uses_stq : _GEN_6965; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_uses_ldq = slots_16_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7164 = _T_905 ? issue_slots_16_uop_uses_ldq : _GEN_6966; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_amo = slots_16_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7165 = _T_905 ? issue_slots_16_uop_is_amo : _GEN_6967; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_fencei = slots_16_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7166 = _T_905 ? issue_slots_16_uop_is_fencei : _GEN_6968; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_fence = slots_16_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7167 = _T_905 ? issue_slots_16_uop_is_fence : _GEN_6969; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_mem_signed = slots_16_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7168 = _T_905 ? issue_slots_16_uop_mem_signed : _GEN_6970; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_mem_size = slots_16_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7169 = _T_905 ? issue_slots_16_uop_mem_size : _GEN_6971; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_16_uop_mem_cmd = slots_16_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7170 = _T_905 ? issue_slots_16_uop_mem_cmd : _GEN_6972; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_bypassable = slots_16_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7171 = _T_905 ? issue_slots_16_uop_bypassable : _GEN_6973; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_16_uop_exc_cause = slots_16_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_7172 = _T_905 ? issue_slots_16_uop_exc_cause : _GEN_6974; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_exception = slots_16_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7173 = _T_905 ? issue_slots_16_uop_exception : _GEN_6975; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_16_uop_stale_pdst = slots_16_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7174 = _T_905 ? issue_slots_16_uop_stale_pdst : _GEN_6976; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_ppred_busy = slots_16_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7175 = _T_905 ? issue_slots_16_uop_ppred_busy : _GEN_6977; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_prs3_busy = slots_16_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7176 = _T_905 ? issue_slots_16_uop_prs3_busy : _GEN_6978; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_prs2_busy = slots_16_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7177 = _T_905 ? issue_slots_16_uop_prs2_busy : _GEN_6979; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_prs1_busy = slots_16_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7178 = _T_905 ? issue_slots_16_uop_prs1_busy : _GEN_6980; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_16_uop_ppred = slots_16_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7179 = _T_905 ? issue_slots_16_uop_ppred : _GEN_6981; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_16_uop_prs3 = slots_16_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7180 = _T_905 ? issue_slots_16_uop_prs3 : _GEN_6982; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_16_uop_prs2 = slots_16_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7181 = _T_905 ? issue_slots_16_uop_prs2 : _GEN_6983; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_16_uop_prs1 = slots_16_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7182 = _T_905 ? issue_slots_16_uop_prs1 : _GEN_6984; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_16_uop_pdst = slots_16_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7183 = _T_905 ? issue_slots_16_uop_pdst : _GEN_6985; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_rxq_idx = slots_16_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7184 = _T_905 ? issue_slots_16_uop_rxq_idx : _GEN_6986; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_16_uop_stq_idx = slots_16_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7185 = _T_905 ? issue_slots_16_uop_stq_idx : _GEN_6987; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_16_uop_ldq_idx = slots_16_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7186 = _T_905 ? issue_slots_16_uop_ldq_idx : _GEN_6988; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_rob_idx = slots_16_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7187 = _T_905 ? issue_slots_16_uop_rob_idx : _GEN_6989; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_16_uop_csr_addr = slots_16_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_7188 = _T_905 ? issue_slots_16_uop_csr_addr : _GEN_6990; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_16_uop_imm_packed = slots_16_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_7189 = _T_905 ? issue_slots_16_uop_imm_packed : _GEN_6991; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_taken = slots_16_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7190 = _T_905 ? issue_slots_16_uop_taken : _GEN_6992; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_pc_lob = slots_16_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7191 = _T_905 ? issue_slots_16_uop_pc_lob : _GEN_6993; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_edge_inst = slots_16_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7192 = _T_905 ? issue_slots_16_uop_edge_inst : _GEN_6994; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_16_uop_ftq_idx = slots_16_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7193 = _T_905 ? issue_slots_16_uop_ftq_idx : _GEN_6995; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_br_tag = slots_16_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7194 = _T_905 ? issue_slots_16_uop_br_tag : _GEN_6996; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_16_uop_br_mask = slots_16_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_7195 = _T_905 ? issue_slots_16_uop_br_mask : _GEN_6997; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_sfb = slots_16_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7196 = _T_905 ? issue_slots_16_uop_is_sfb : _GEN_6998; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_jal = slots_16_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7197 = _T_905 ? issue_slots_16_uop_is_jal : _GEN_6999; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_jalr = slots_16_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7198 = _T_905 ? issue_slots_16_uop_is_jalr : _GEN_7000; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_br = slots_16_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7199 = _T_905 ? issue_slots_16_uop_is_br : _GEN_7001; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_iw_p2_poisoned = slots_16_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7200 = _T_905 ? issue_slots_16_uop_iw_p2_poisoned : _GEN_7002; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_iw_p1_poisoned = slots_16_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7201 = _T_905 ? issue_slots_16_uop_iw_p1_poisoned : _GEN_7003; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_iw_state = slots_16_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7202 = _T_905 ? issue_slots_16_uop_iw_state : _GEN_7004; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_ctrl_op3_sel = slots_16_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7203 = _T_905 ? issue_slots_16_uop_ctrl_op3_sel : _GEN_7005; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_ctrl_is_std = slots_16_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7204 = _T_905 ? issue_slots_16_uop_ctrl_is_std : _GEN_7006; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_ctrl_is_sta = slots_16_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7205 = _T_905 ? issue_slots_16_uop_ctrl_is_sta : _GEN_7007; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_ctrl_is_load = slots_16_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7206 = _T_905 ? issue_slots_16_uop_ctrl_is_load : _GEN_7008; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_16_uop_ctrl_csr_cmd = slots_16_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7207 = _T_905 ? issue_slots_16_uop_ctrl_csr_cmd : _GEN_7009; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_ctrl_fcn_dw = slots_16_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7208 = _T_905 ? issue_slots_16_uop_ctrl_fcn_dw : _GEN_7010; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_ctrl_op_fcn = slots_16_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7209 = _T_905 ? issue_slots_16_uop_ctrl_op_fcn : _GEN_7011; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_16_uop_ctrl_imm_sel = slots_16_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7210 = _T_905 ? issue_slots_16_uop_ctrl_imm_sel : _GEN_7012; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_16_uop_ctrl_op2_sel = slots_16_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7211 = _T_905 ? issue_slots_16_uop_ctrl_op2_sel : _GEN_7013; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_ctrl_op1_sel = slots_16_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7212 = _T_905 ? issue_slots_16_uop_ctrl_op1_sel : _GEN_7014; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_ctrl_br_type = slots_16_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7213 = _T_905 ? issue_slots_16_uop_ctrl_br_type : _GEN_7015; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7214 = _T_905 ? issue_slots_16_uop_fu_code : _GEN_7016; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_16_uop_iq_type = slots_16_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7215 = _T_905 ? issue_slots_16_uop_iq_type : _GEN_7017; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_16_uop_debug_pc = slots_16_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_7216 = _T_905 ? issue_slots_16_uop_debug_pc : _GEN_7018; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_rvc = slots_16_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7217 = _T_905 ? issue_slots_16_uop_is_rvc : _GEN_7019; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_16_uop_debug_inst = slots_16_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7218 = _T_905 ? issue_slots_16_uop_debug_inst : _GEN_7020; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_16_uop_inst = slots_16_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7219 = _T_905 ? issue_slots_16_uop_inst : _GEN_7021; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_16_uop_uopc = slots_16_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7220 = _T_905 ? issue_slots_16_uop_uopc : _GEN_7022; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_address_num = slots_16_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7221 = _T_905 ? issue_slots_16_uop_address_num : _GEN_7023; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_rob_inst_idx = slots_16_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7222 = _T_905 ? issue_slots_16_uop_rob_inst_idx : _GEN_7024; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_self_index = slots_16_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7223 = _T_905 ? issue_slots_16_uop_self_index : _GEN_7025; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_16_uop_split_num = slots_16_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7224 = _T_905 ? issue_slots_16_uop_split_num : _GEN_7026; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_op2_sel = slots_16_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7225 = _T_905 ? issue_slots_16_uop_op2_sel : _GEN_7027; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_op1_sel = slots_16_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7226 = _T_905 ? issue_slots_16_uop_op1_sel : _GEN_7028; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_stale_pflag = slots_16_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7227 = _T_905 ? issue_slots_16_uop_stale_pflag : _GEN_7029; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_pflag_busy = slots_16_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7228 = _T_905 ? issue_slots_16_uop_pflag_busy : _GEN_7030; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_pwflag = slots_16_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7229 = _T_905 ? issue_slots_16_uop_pwflag : _GEN_7031; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_16_uop_prflag = slots_16_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7230 = _T_905 ? issue_slots_16_uop_prflag : _GEN_7032; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_wflag = slots_16_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7231 = _T_905 ? issue_slots_16_uop_wflag : _GEN_7033; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_rflag = slots_16_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7232 = _T_905 ? issue_slots_16_uop_rflag : _GEN_7034; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_16_uop_lrs3_rtype = slots_16_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7233 = _T_905 ? issue_slots_16_uop_lrs3_rtype : _GEN_7035; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_16_uop_shift = slots_16_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7234 = _T_905 ? issue_slots_16_uop_shift : _GEN_7036; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_is_unicore = slots_16_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7235 = _T_905 ? issue_slots_16_uop_is_unicore : _GEN_7037; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_switch_off = slots_16_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7236 = _T_905 ? issue_slots_16_uop_switch_off : _GEN_7038; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_16_uop_switch = slots_16_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7237 = _T_905 ? issue_slots_16_uop_switch : _GEN_7039; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7240 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_debug_tsrc : _GEN_7042
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7241 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_debug_fsrc : _GEN_7043
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7242 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_bp_xcpt_if : _GEN_7044; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7243 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_bp_debug_if : _GEN_7045; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7244 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_xcpt_ma_if : _GEN_7046; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7245 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_xcpt_ae_if : _GEN_7047; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7246 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_xcpt_pf_if : _GEN_7048; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7247 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_fp_single : _GEN_7049; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7248 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_fp_val : _GEN_7050; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7249 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_frs3_en : _GEN_7051; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7250 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_lrs2_rtype : _GEN_7052
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7251 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_lrs1_rtype : _GEN_7053
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7252 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_dst_rtype : _GEN_7054; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7253 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ldst_val : _GEN_7055; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7254 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_lrs3 : _GEN_7056; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7255 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_lrs2 : _GEN_7057; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7256 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_lrs1 : _GEN_7058; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7257 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ldst : _GEN_7059; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7258 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ldst_is_rs1 : _GEN_7060; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7259 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_flush_on_commit : _GEN_7061
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7260 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_unique : _GEN_7062; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7261 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_sys_pc2epc : _GEN_7063; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7262 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_uses_stq : _GEN_7064; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7263 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_uses_ldq : _GEN_7065; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7264 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_amo : _GEN_7066; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7265 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_fencei : _GEN_7067; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7266 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_fence : _GEN_7068; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7267 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_mem_signed : _GEN_7069; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7268 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_mem_size : _GEN_7070; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7269 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_mem_cmd : _GEN_7071; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7270 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_bypassable : _GEN_7072; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_7271 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_exc_cause : _GEN_7073
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7272 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_exception : _GEN_7074; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7273 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_stale_pdst : _GEN_7075
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7274 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ppred_busy : _GEN_7076; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7275 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_prs3_busy : _GEN_7077; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7276 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_prs2_busy : _GEN_7078; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7277 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_prs1_busy : _GEN_7079; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7278 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ppred : _GEN_7080; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7279 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_prs3 : _GEN_7081; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7280 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_prs2 : _GEN_7082; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7281 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_prs1 : _GEN_7083; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7282 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_pdst : _GEN_7084; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7283 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_rxq_idx : _GEN_7085; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7284 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_stq_idx : _GEN_7086; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7285 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ldq_idx : _GEN_7087; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7286 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_rob_idx : _GEN_7088; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7287 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_csr_addr : _GEN_7089; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_7288 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_imm_packed :
    _GEN_7090; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7289 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_taken : _GEN_7091; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7290 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_pc_lob : _GEN_7092; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7291 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_edge_inst : _GEN_7093; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7292 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ftq_idx : _GEN_7094; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7293 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_br_tag : _GEN_7095; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7294 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_br_mask : _GEN_7096; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7295 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_sfb : _GEN_7097; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7296 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_jal : _GEN_7098; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7297 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_jalr : _GEN_7099; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7298 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_br : _GEN_7100; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7299 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_iw_p2_poisoned : _GEN_7101; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7300 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_iw_p1_poisoned : _GEN_7102; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7301 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_iw_state : _GEN_7103; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7302 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_op3_sel :
    _GEN_7104; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7303 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_is_std : _GEN_7105; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7304 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_is_sta : _GEN_7106; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7305 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_is_load : _GEN_7107; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7306 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_csr_cmd :
    _GEN_7108; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7307 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_fcn_dw : _GEN_7109; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7308 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_op_fcn :
    _GEN_7110; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7309 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_imm_sel :
    _GEN_7111; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7310 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_op2_sel :
    _GEN_7112; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7311 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_op1_sel :
    _GEN_7113; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7312 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_ctrl_br_type :
    _GEN_7114; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7313 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_fu_code : _GEN_7115; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7314 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_iq_type : _GEN_7116; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_7315 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_debug_pc : _GEN_7117; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7316 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_rvc : _GEN_7118; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7317 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_debug_inst :
    _GEN_7119; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7318 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_inst : _GEN_7120; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7319 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_uopc : _GEN_7121; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7320 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_address_num :
    _GEN_7122; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7321 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_rob_inst_idx :
    _GEN_7123; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7322 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_self_index : _GEN_7124
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7323 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_split_num : _GEN_7125; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7324 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_op2_sel : _GEN_7126; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7325 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_op1_sel : _GEN_7127; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7326 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_stale_pflag :
    _GEN_7128; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7327 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_pflag_busy : _GEN_7129; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7328 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_pwflag : _GEN_7130; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7329 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_prflag : _GEN_7131; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7330 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_wflag : _GEN_7132; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7331 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_rflag : _GEN_7133; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7332 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_lrs3_rtype : _GEN_7134
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7333 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_shift : _GEN_7135; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7334 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_is_unicore : _GEN_7136; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7335 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_switch_off : _GEN_7137; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7336 = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 ? issue_slots_16_uop_switch : _GEN_7138; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_debug_tsrc = slots_17_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7339 = _T_935 ? issue_slots_17_uop_debug_tsrc : _GEN_7141; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_debug_fsrc = slots_17_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7340 = _T_935 ? issue_slots_17_uop_debug_fsrc : _GEN_7142; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_bp_xcpt_if = slots_17_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7341 = _T_935 ? issue_slots_17_uop_bp_xcpt_if : _GEN_7143; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_bp_debug_if = slots_17_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7342 = _T_935 ? issue_slots_17_uop_bp_debug_if : _GEN_7144; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_xcpt_ma_if = slots_17_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7343 = _T_935 ? issue_slots_17_uop_xcpt_ma_if : _GEN_7145; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_xcpt_ae_if = slots_17_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7344 = _T_935 ? issue_slots_17_uop_xcpt_ae_if : _GEN_7146; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_xcpt_pf_if = slots_17_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7345 = _T_935 ? issue_slots_17_uop_xcpt_pf_if : _GEN_7147; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_fp_single = slots_17_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7346 = _T_935 ? issue_slots_17_uop_fp_single : _GEN_7148; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_fp_val = slots_17_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7347 = _T_935 ? issue_slots_17_uop_fp_val : _GEN_7149; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_frs3_en = slots_17_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7348 = _T_935 ? issue_slots_17_uop_frs3_en : _GEN_7150; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_lrs2_rtype = slots_17_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7349 = _T_935 ? issue_slots_17_uop_lrs2_rtype : _GEN_7151; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_lrs1_rtype = slots_17_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7350 = _T_935 ? issue_slots_17_uop_lrs1_rtype : _GEN_7152; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_dst_rtype = slots_17_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7351 = _T_935 ? issue_slots_17_uop_dst_rtype : _GEN_7153; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_ldst_val = slots_17_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7352 = _T_935 ? issue_slots_17_uop_ldst_val : _GEN_7154; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_lrs3 = slots_17_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7353 = _T_935 ? issue_slots_17_uop_lrs3 : _GEN_7155; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_lrs2 = slots_17_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7354 = _T_935 ? issue_slots_17_uop_lrs2 : _GEN_7156; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_lrs1 = slots_17_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7355 = _T_935 ? issue_slots_17_uop_lrs1 : _GEN_7157; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_ldst = slots_17_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7356 = _T_935 ? issue_slots_17_uop_ldst : _GEN_7158; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_ldst_is_rs1 = slots_17_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7357 = _T_935 ? issue_slots_17_uop_ldst_is_rs1 : _GEN_7159; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_flush_on_commit = slots_17_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7358 = _T_935 ? issue_slots_17_uop_flush_on_commit : _GEN_7160; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_unique = slots_17_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7359 = _T_935 ? issue_slots_17_uop_is_unique : _GEN_7161; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_sys_pc2epc = slots_17_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7360 = _T_935 ? issue_slots_17_uop_is_sys_pc2epc : _GEN_7162; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_uses_stq = slots_17_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7361 = _T_935 ? issue_slots_17_uop_uses_stq : _GEN_7163; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_uses_ldq = slots_17_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7362 = _T_935 ? issue_slots_17_uop_uses_ldq : _GEN_7164; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_amo = slots_17_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7363 = _T_935 ? issue_slots_17_uop_is_amo : _GEN_7165; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_fencei = slots_17_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7364 = _T_935 ? issue_slots_17_uop_is_fencei : _GEN_7166; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_fence = slots_17_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7365 = _T_935 ? issue_slots_17_uop_is_fence : _GEN_7167; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_mem_signed = slots_17_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7366 = _T_935 ? issue_slots_17_uop_mem_signed : _GEN_7168; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_mem_size = slots_17_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7367 = _T_935 ? issue_slots_17_uop_mem_size : _GEN_7169; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_17_uop_mem_cmd = slots_17_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7368 = _T_935 ? issue_slots_17_uop_mem_cmd : _GEN_7170; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_bypassable = slots_17_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7369 = _T_935 ? issue_slots_17_uop_bypassable : _GEN_7171; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_17_uop_exc_cause = slots_17_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_7370 = _T_935 ? issue_slots_17_uop_exc_cause : _GEN_7172; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_exception = slots_17_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7371 = _T_935 ? issue_slots_17_uop_exception : _GEN_7173; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_17_uop_stale_pdst = slots_17_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7372 = _T_935 ? issue_slots_17_uop_stale_pdst : _GEN_7174; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_ppred_busy = slots_17_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7373 = _T_935 ? issue_slots_17_uop_ppred_busy : _GEN_7175; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_prs3_busy = slots_17_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7374 = _T_935 ? issue_slots_17_uop_prs3_busy : _GEN_7176; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_prs2_busy = slots_17_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7375 = _T_935 ? issue_slots_17_uop_prs2_busy : _GEN_7177; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_prs1_busy = slots_17_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7376 = _T_935 ? issue_slots_17_uop_prs1_busy : _GEN_7178; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_17_uop_ppred = slots_17_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7377 = _T_935 ? issue_slots_17_uop_ppred : _GEN_7179; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_17_uop_prs3 = slots_17_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7378 = _T_935 ? issue_slots_17_uop_prs3 : _GEN_7180; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_17_uop_prs2 = slots_17_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7379 = _T_935 ? issue_slots_17_uop_prs2 : _GEN_7181; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_17_uop_prs1 = slots_17_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7380 = _T_935 ? issue_slots_17_uop_prs1 : _GEN_7182; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_17_uop_pdst = slots_17_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7381 = _T_935 ? issue_slots_17_uop_pdst : _GEN_7183; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_rxq_idx = slots_17_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7382 = _T_935 ? issue_slots_17_uop_rxq_idx : _GEN_7184; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_17_uop_stq_idx = slots_17_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7383 = _T_935 ? issue_slots_17_uop_stq_idx : _GEN_7185; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_17_uop_ldq_idx = slots_17_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7384 = _T_935 ? issue_slots_17_uop_ldq_idx : _GEN_7186; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_rob_idx = slots_17_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7385 = _T_935 ? issue_slots_17_uop_rob_idx : _GEN_7187; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_17_uop_csr_addr = slots_17_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_7386 = _T_935 ? issue_slots_17_uop_csr_addr : _GEN_7188; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_17_uop_imm_packed = slots_17_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_7387 = _T_935 ? issue_slots_17_uop_imm_packed : _GEN_7189; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_taken = slots_17_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7388 = _T_935 ? issue_slots_17_uop_taken : _GEN_7190; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_pc_lob = slots_17_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7389 = _T_935 ? issue_slots_17_uop_pc_lob : _GEN_7191; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_edge_inst = slots_17_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7390 = _T_935 ? issue_slots_17_uop_edge_inst : _GEN_7192; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_17_uop_ftq_idx = slots_17_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7391 = _T_935 ? issue_slots_17_uop_ftq_idx : _GEN_7193; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_br_tag = slots_17_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7392 = _T_935 ? issue_slots_17_uop_br_tag : _GEN_7194; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_17_uop_br_mask = slots_17_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_7393 = _T_935 ? issue_slots_17_uop_br_mask : _GEN_7195; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_sfb = slots_17_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7394 = _T_935 ? issue_slots_17_uop_is_sfb : _GEN_7196; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_jal = slots_17_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7395 = _T_935 ? issue_slots_17_uop_is_jal : _GEN_7197; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_jalr = slots_17_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7396 = _T_935 ? issue_slots_17_uop_is_jalr : _GEN_7198; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_br = slots_17_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7397 = _T_935 ? issue_slots_17_uop_is_br : _GEN_7199; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_iw_p2_poisoned = slots_17_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7398 = _T_935 ? issue_slots_17_uop_iw_p2_poisoned : _GEN_7200; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_iw_p1_poisoned = slots_17_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7399 = _T_935 ? issue_slots_17_uop_iw_p1_poisoned : _GEN_7201; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_iw_state = slots_17_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7400 = _T_935 ? issue_slots_17_uop_iw_state : _GEN_7202; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_ctrl_op3_sel = slots_17_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7401 = _T_935 ? issue_slots_17_uop_ctrl_op3_sel : _GEN_7203; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_ctrl_is_std = slots_17_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7402 = _T_935 ? issue_slots_17_uop_ctrl_is_std : _GEN_7204; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_ctrl_is_sta = slots_17_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7403 = _T_935 ? issue_slots_17_uop_ctrl_is_sta : _GEN_7205; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_ctrl_is_load = slots_17_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7404 = _T_935 ? issue_slots_17_uop_ctrl_is_load : _GEN_7206; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_17_uop_ctrl_csr_cmd = slots_17_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7405 = _T_935 ? issue_slots_17_uop_ctrl_csr_cmd : _GEN_7207; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_ctrl_fcn_dw = slots_17_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7406 = _T_935 ? issue_slots_17_uop_ctrl_fcn_dw : _GEN_7208; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_ctrl_op_fcn = slots_17_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7407 = _T_935 ? issue_slots_17_uop_ctrl_op_fcn : _GEN_7209; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_17_uop_ctrl_imm_sel = slots_17_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7408 = _T_935 ? issue_slots_17_uop_ctrl_imm_sel : _GEN_7210; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_17_uop_ctrl_op2_sel = slots_17_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7409 = _T_935 ? issue_slots_17_uop_ctrl_op2_sel : _GEN_7211; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_ctrl_op1_sel = slots_17_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7410 = _T_935 ? issue_slots_17_uop_ctrl_op1_sel : _GEN_7212; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_ctrl_br_type = slots_17_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7411 = _T_935 ? issue_slots_17_uop_ctrl_br_type : _GEN_7213; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7412 = _T_935 ? issue_slots_17_uop_fu_code : _GEN_7214; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_17_uop_iq_type = slots_17_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7413 = _T_935 ? issue_slots_17_uop_iq_type : _GEN_7215; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_17_uop_debug_pc = slots_17_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_7414 = _T_935 ? issue_slots_17_uop_debug_pc : _GEN_7216; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_rvc = slots_17_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7415 = _T_935 ? issue_slots_17_uop_is_rvc : _GEN_7217; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_17_uop_debug_inst = slots_17_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7416 = _T_935 ? issue_slots_17_uop_debug_inst : _GEN_7218; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_17_uop_inst = slots_17_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7417 = _T_935 ? issue_slots_17_uop_inst : _GEN_7219; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_17_uop_uopc = slots_17_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7418 = _T_935 ? issue_slots_17_uop_uopc : _GEN_7220; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_address_num = slots_17_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7419 = _T_935 ? issue_slots_17_uop_address_num : _GEN_7221; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_rob_inst_idx = slots_17_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7420 = _T_935 ? issue_slots_17_uop_rob_inst_idx : _GEN_7222; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_self_index = slots_17_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7421 = _T_935 ? issue_slots_17_uop_self_index : _GEN_7223; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_17_uop_split_num = slots_17_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7422 = _T_935 ? issue_slots_17_uop_split_num : _GEN_7224; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_op2_sel = slots_17_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7423 = _T_935 ? issue_slots_17_uop_op2_sel : _GEN_7225; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_op1_sel = slots_17_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7424 = _T_935 ? issue_slots_17_uop_op1_sel : _GEN_7226; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_stale_pflag = slots_17_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7425 = _T_935 ? issue_slots_17_uop_stale_pflag : _GEN_7227; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_pflag_busy = slots_17_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7426 = _T_935 ? issue_slots_17_uop_pflag_busy : _GEN_7228; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_pwflag = slots_17_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7427 = _T_935 ? issue_slots_17_uop_pwflag : _GEN_7229; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_17_uop_prflag = slots_17_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7428 = _T_935 ? issue_slots_17_uop_prflag : _GEN_7230; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_wflag = slots_17_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7429 = _T_935 ? issue_slots_17_uop_wflag : _GEN_7231; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_rflag = slots_17_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7430 = _T_935 ? issue_slots_17_uop_rflag : _GEN_7232; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_17_uop_lrs3_rtype = slots_17_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7431 = _T_935 ? issue_slots_17_uop_lrs3_rtype : _GEN_7233; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_17_uop_shift = slots_17_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7432 = _T_935 ? issue_slots_17_uop_shift : _GEN_7234; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_is_unicore = slots_17_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7433 = _T_935 ? issue_slots_17_uop_is_unicore : _GEN_7235; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_switch_off = slots_17_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7434 = _T_935 ? issue_slots_17_uop_switch_off : _GEN_7236; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_17_uop_switch = slots_17_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7435 = _T_935 ? issue_slots_17_uop_switch : _GEN_7237; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7438 = _T_946 & ~_T_917 ? issue_slots_17_uop_debug_tsrc : _GEN_7240; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7439 = _T_946 & ~_T_917 ? issue_slots_17_uop_debug_fsrc : _GEN_7241; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7440 = _T_946 & ~_T_917 ? issue_slots_17_uop_bp_xcpt_if : _GEN_7242; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7441 = _T_946 & ~_T_917 ? issue_slots_17_uop_bp_debug_if : _GEN_7243; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7442 = _T_946 & ~_T_917 ? issue_slots_17_uop_xcpt_ma_if : _GEN_7244; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7443 = _T_946 & ~_T_917 ? issue_slots_17_uop_xcpt_ae_if : _GEN_7245; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7444 = _T_946 & ~_T_917 ? issue_slots_17_uop_xcpt_pf_if : _GEN_7246; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7445 = _T_946 & ~_T_917 ? issue_slots_17_uop_fp_single : _GEN_7247; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7446 = _T_946 & ~_T_917 ? issue_slots_17_uop_fp_val : _GEN_7248; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7447 = _T_946 & ~_T_917 ? issue_slots_17_uop_frs3_en : _GEN_7249; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7448 = _T_946 & ~_T_917 ? issue_slots_17_uop_lrs2_rtype : _GEN_7250; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7449 = _T_946 & ~_T_917 ? issue_slots_17_uop_lrs1_rtype : _GEN_7251; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7450 = _T_946 & ~_T_917 ? issue_slots_17_uop_dst_rtype : _GEN_7252; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7451 = _T_946 & ~_T_917 ? issue_slots_17_uop_ldst_val : _GEN_7253; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7452 = _T_946 & ~_T_917 ? issue_slots_17_uop_lrs3 : _GEN_7254; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7453 = _T_946 & ~_T_917 ? issue_slots_17_uop_lrs2 : _GEN_7255; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7454 = _T_946 & ~_T_917 ? issue_slots_17_uop_lrs1 : _GEN_7256; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7455 = _T_946 & ~_T_917 ? issue_slots_17_uop_ldst : _GEN_7257; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7456 = _T_946 & ~_T_917 ? issue_slots_17_uop_ldst_is_rs1 : _GEN_7258; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7457 = _T_946 & ~_T_917 ? issue_slots_17_uop_flush_on_commit : _GEN_7259; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7458 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_unique : _GEN_7260; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7459 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_sys_pc2epc : _GEN_7261; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7460 = _T_946 & ~_T_917 ? issue_slots_17_uop_uses_stq : _GEN_7262; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7461 = _T_946 & ~_T_917 ? issue_slots_17_uop_uses_ldq : _GEN_7263; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7462 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_amo : _GEN_7264; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7463 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_fencei : _GEN_7265; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7464 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_fence : _GEN_7266; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7465 = _T_946 & ~_T_917 ? issue_slots_17_uop_mem_signed : _GEN_7267; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7466 = _T_946 & ~_T_917 ? issue_slots_17_uop_mem_size : _GEN_7268; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7467 = _T_946 & ~_T_917 ? issue_slots_17_uop_mem_cmd : _GEN_7269; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7468 = _T_946 & ~_T_917 ? issue_slots_17_uop_bypassable : _GEN_7270; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_7469 = _T_946 & ~_T_917 ? issue_slots_17_uop_exc_cause : _GEN_7271; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7470 = _T_946 & ~_T_917 ? issue_slots_17_uop_exception : _GEN_7272; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7471 = _T_946 & ~_T_917 ? issue_slots_17_uop_stale_pdst : _GEN_7273; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7472 = _T_946 & ~_T_917 ? issue_slots_17_uop_ppred_busy : _GEN_7274; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7473 = _T_946 & ~_T_917 ? issue_slots_17_uop_prs3_busy : _GEN_7275; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7474 = _T_946 & ~_T_917 ? issue_slots_17_uop_prs2_busy : _GEN_7276; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7475 = _T_946 & ~_T_917 ? issue_slots_17_uop_prs1_busy : _GEN_7277; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7476 = _T_946 & ~_T_917 ? issue_slots_17_uop_ppred : _GEN_7278; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7477 = _T_946 & ~_T_917 ? issue_slots_17_uop_prs3 : _GEN_7279; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7478 = _T_946 & ~_T_917 ? issue_slots_17_uop_prs2 : _GEN_7280; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7479 = _T_946 & ~_T_917 ? issue_slots_17_uop_prs1 : _GEN_7281; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7480 = _T_946 & ~_T_917 ? issue_slots_17_uop_pdst : _GEN_7282; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7481 = _T_946 & ~_T_917 ? issue_slots_17_uop_rxq_idx : _GEN_7283; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7482 = _T_946 & ~_T_917 ? issue_slots_17_uop_stq_idx : _GEN_7284; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7483 = _T_946 & ~_T_917 ? issue_slots_17_uop_ldq_idx : _GEN_7285; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7484 = _T_946 & ~_T_917 ? issue_slots_17_uop_rob_idx : _GEN_7286; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7485 = _T_946 & ~_T_917 ? issue_slots_17_uop_csr_addr : _GEN_7287; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_7486 = _T_946 & ~_T_917 ? issue_slots_17_uop_imm_packed : _GEN_7288; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7487 = _T_946 & ~_T_917 ? issue_slots_17_uop_taken : _GEN_7289; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7488 = _T_946 & ~_T_917 ? issue_slots_17_uop_pc_lob : _GEN_7290; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7489 = _T_946 & ~_T_917 ? issue_slots_17_uop_edge_inst : _GEN_7291; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7490 = _T_946 & ~_T_917 ? issue_slots_17_uop_ftq_idx : _GEN_7292; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7491 = _T_946 & ~_T_917 ? issue_slots_17_uop_br_tag : _GEN_7293; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7492 = _T_946 & ~_T_917 ? issue_slots_17_uop_br_mask : _GEN_7294; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7493 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_sfb : _GEN_7295; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7494 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_jal : _GEN_7296; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7495 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_jalr : _GEN_7297; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7496 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_br : _GEN_7298; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7497 = _T_946 & ~_T_917 ? issue_slots_17_uop_iw_p2_poisoned : _GEN_7299; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7498 = _T_946 & ~_T_917 ? issue_slots_17_uop_iw_p1_poisoned : _GEN_7300; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7499 = _T_946 & ~_T_917 ? issue_slots_17_uop_iw_state : _GEN_7301; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7500 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_op3_sel : _GEN_7302; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7501 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_is_std : _GEN_7303; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7502 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_is_sta : _GEN_7304; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7503 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_is_load : _GEN_7305; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7504 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_csr_cmd : _GEN_7306; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7505 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_fcn_dw : _GEN_7307; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7506 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_op_fcn : _GEN_7308; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7507 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_imm_sel : _GEN_7309; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7508 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_op2_sel : _GEN_7310; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7509 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_op1_sel : _GEN_7311; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7510 = _T_946 & ~_T_917 ? issue_slots_17_uop_ctrl_br_type : _GEN_7312; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7511 = _T_946 & ~_T_917 ? issue_slots_17_uop_fu_code : _GEN_7313; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7512 = _T_946 & ~_T_917 ? issue_slots_17_uop_iq_type : _GEN_7314; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_7513 = _T_946 & ~_T_917 ? issue_slots_17_uop_debug_pc : _GEN_7315; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7514 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_rvc : _GEN_7316; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7515 = _T_946 & ~_T_917 ? issue_slots_17_uop_debug_inst : _GEN_7317; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7516 = _T_946 & ~_T_917 ? issue_slots_17_uop_inst : _GEN_7318; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7517 = _T_946 & ~_T_917 ? issue_slots_17_uop_uopc : _GEN_7319; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7518 = _T_946 & ~_T_917 ? issue_slots_17_uop_address_num : _GEN_7320; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7519 = _T_946 & ~_T_917 ? issue_slots_17_uop_rob_inst_idx : _GEN_7321; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7520 = _T_946 & ~_T_917 ? issue_slots_17_uop_self_index : _GEN_7322; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7521 = _T_946 & ~_T_917 ? issue_slots_17_uop_split_num : _GEN_7323; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7522 = _T_946 & ~_T_917 ? issue_slots_17_uop_op2_sel : _GEN_7324; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7523 = _T_946 & ~_T_917 ? issue_slots_17_uop_op1_sel : _GEN_7325; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7524 = _T_946 & ~_T_917 ? issue_slots_17_uop_stale_pflag : _GEN_7326; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7525 = _T_946 & ~_T_917 ? issue_slots_17_uop_pflag_busy : _GEN_7327; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7526 = _T_946 & ~_T_917 ? issue_slots_17_uop_pwflag : _GEN_7328; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7527 = _T_946 & ~_T_917 ? issue_slots_17_uop_prflag : _GEN_7329; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7528 = _T_946 & ~_T_917 ? issue_slots_17_uop_wflag : _GEN_7330; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7529 = _T_946 & ~_T_917 ? issue_slots_17_uop_rflag : _GEN_7331; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7530 = _T_946 & ~_T_917 ? issue_slots_17_uop_lrs3_rtype : _GEN_7332; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7531 = _T_946 & ~_T_917 ? issue_slots_17_uop_shift : _GEN_7333; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7532 = _T_946 & ~_T_917 ? issue_slots_17_uop_is_unicore : _GEN_7334; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7533 = _T_946 & ~_T_917 ? issue_slots_17_uop_switch_off : _GEN_7335; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7534 = _T_946 & ~_T_917 ? issue_slots_17_uop_switch : _GEN_7336; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_debug_tsrc = slots_18_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7537 = _T_965 ? issue_slots_18_uop_debug_tsrc : _GEN_7339; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_debug_fsrc = slots_18_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7538 = _T_965 ? issue_slots_18_uop_debug_fsrc : _GEN_7340; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_bp_xcpt_if = slots_18_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7539 = _T_965 ? issue_slots_18_uop_bp_xcpt_if : _GEN_7341; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_bp_debug_if = slots_18_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7540 = _T_965 ? issue_slots_18_uop_bp_debug_if : _GEN_7342; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_xcpt_ma_if = slots_18_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7541 = _T_965 ? issue_slots_18_uop_xcpt_ma_if : _GEN_7343; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_xcpt_ae_if = slots_18_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7542 = _T_965 ? issue_slots_18_uop_xcpt_ae_if : _GEN_7344; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_xcpt_pf_if = slots_18_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7543 = _T_965 ? issue_slots_18_uop_xcpt_pf_if : _GEN_7345; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_fp_single = slots_18_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7544 = _T_965 ? issue_slots_18_uop_fp_single : _GEN_7346; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_fp_val = slots_18_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7545 = _T_965 ? issue_slots_18_uop_fp_val : _GEN_7347; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_frs3_en = slots_18_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7546 = _T_965 ? issue_slots_18_uop_frs3_en : _GEN_7348; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_lrs2_rtype = slots_18_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7547 = _T_965 ? issue_slots_18_uop_lrs2_rtype : _GEN_7349; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_lrs1_rtype = slots_18_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7548 = _T_965 ? issue_slots_18_uop_lrs1_rtype : _GEN_7350; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_dst_rtype = slots_18_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7549 = _T_965 ? issue_slots_18_uop_dst_rtype : _GEN_7351; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_ldst_val = slots_18_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7550 = _T_965 ? issue_slots_18_uop_ldst_val : _GEN_7352; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_lrs3 = slots_18_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7551 = _T_965 ? issue_slots_18_uop_lrs3 : _GEN_7353; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_lrs2 = slots_18_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7552 = _T_965 ? issue_slots_18_uop_lrs2 : _GEN_7354; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_lrs1 = slots_18_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7553 = _T_965 ? issue_slots_18_uop_lrs1 : _GEN_7355; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_ldst = slots_18_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7554 = _T_965 ? issue_slots_18_uop_ldst : _GEN_7356; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_ldst_is_rs1 = slots_18_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7555 = _T_965 ? issue_slots_18_uop_ldst_is_rs1 : _GEN_7357; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_flush_on_commit = slots_18_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7556 = _T_965 ? issue_slots_18_uop_flush_on_commit : _GEN_7358; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_unique = slots_18_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7557 = _T_965 ? issue_slots_18_uop_is_unique : _GEN_7359; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_sys_pc2epc = slots_18_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7558 = _T_965 ? issue_slots_18_uop_is_sys_pc2epc : _GEN_7360; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_uses_stq = slots_18_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7559 = _T_965 ? issue_slots_18_uop_uses_stq : _GEN_7361; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_uses_ldq = slots_18_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7560 = _T_965 ? issue_slots_18_uop_uses_ldq : _GEN_7362; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_amo = slots_18_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7561 = _T_965 ? issue_slots_18_uop_is_amo : _GEN_7363; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_fencei = slots_18_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7562 = _T_965 ? issue_slots_18_uop_is_fencei : _GEN_7364; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_fence = slots_18_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7563 = _T_965 ? issue_slots_18_uop_is_fence : _GEN_7365; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_mem_signed = slots_18_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7564 = _T_965 ? issue_slots_18_uop_mem_signed : _GEN_7366; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_mem_size = slots_18_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7565 = _T_965 ? issue_slots_18_uop_mem_size : _GEN_7367; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_18_uop_mem_cmd = slots_18_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7566 = _T_965 ? issue_slots_18_uop_mem_cmd : _GEN_7368; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_bypassable = slots_18_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7567 = _T_965 ? issue_slots_18_uop_bypassable : _GEN_7369; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_18_uop_exc_cause = slots_18_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_7568 = _T_965 ? issue_slots_18_uop_exc_cause : _GEN_7370; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_exception = slots_18_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7569 = _T_965 ? issue_slots_18_uop_exception : _GEN_7371; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_18_uop_stale_pdst = slots_18_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7570 = _T_965 ? issue_slots_18_uop_stale_pdst : _GEN_7372; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_ppred_busy = slots_18_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7571 = _T_965 ? issue_slots_18_uop_ppred_busy : _GEN_7373; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_prs3_busy = slots_18_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7572 = _T_965 ? issue_slots_18_uop_prs3_busy : _GEN_7374; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_prs2_busy = slots_18_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7573 = _T_965 ? issue_slots_18_uop_prs2_busy : _GEN_7375; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_prs1_busy = slots_18_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7574 = _T_965 ? issue_slots_18_uop_prs1_busy : _GEN_7376; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_18_uop_ppred = slots_18_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7575 = _T_965 ? issue_slots_18_uop_ppred : _GEN_7377; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_18_uop_prs3 = slots_18_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7576 = _T_965 ? issue_slots_18_uop_prs3 : _GEN_7378; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_18_uop_prs2 = slots_18_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7577 = _T_965 ? issue_slots_18_uop_prs2 : _GEN_7379; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_18_uop_prs1 = slots_18_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7578 = _T_965 ? issue_slots_18_uop_prs1 : _GEN_7380; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_18_uop_pdst = slots_18_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7579 = _T_965 ? issue_slots_18_uop_pdst : _GEN_7381; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_rxq_idx = slots_18_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7580 = _T_965 ? issue_slots_18_uop_rxq_idx : _GEN_7382; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_18_uop_stq_idx = slots_18_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7581 = _T_965 ? issue_slots_18_uop_stq_idx : _GEN_7383; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_18_uop_ldq_idx = slots_18_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7582 = _T_965 ? issue_slots_18_uop_ldq_idx : _GEN_7384; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_rob_idx = slots_18_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7583 = _T_965 ? issue_slots_18_uop_rob_idx : _GEN_7385; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_18_uop_csr_addr = slots_18_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_7584 = _T_965 ? issue_slots_18_uop_csr_addr : _GEN_7386; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_18_uop_imm_packed = slots_18_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_7585 = _T_965 ? issue_slots_18_uop_imm_packed : _GEN_7387; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_taken = slots_18_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7586 = _T_965 ? issue_slots_18_uop_taken : _GEN_7388; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_pc_lob = slots_18_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7587 = _T_965 ? issue_slots_18_uop_pc_lob : _GEN_7389; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_edge_inst = slots_18_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7588 = _T_965 ? issue_slots_18_uop_edge_inst : _GEN_7390; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_18_uop_ftq_idx = slots_18_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_7589 = _T_965 ? issue_slots_18_uop_ftq_idx : _GEN_7391; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_br_tag = slots_18_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7590 = _T_965 ? issue_slots_18_uop_br_tag : _GEN_7392; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_18_uop_br_mask = slots_18_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_7591 = _T_965 ? issue_slots_18_uop_br_mask : _GEN_7393; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_sfb = slots_18_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7592 = _T_965 ? issue_slots_18_uop_is_sfb : _GEN_7394; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_jal = slots_18_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7593 = _T_965 ? issue_slots_18_uop_is_jal : _GEN_7395; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_jalr = slots_18_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7594 = _T_965 ? issue_slots_18_uop_is_jalr : _GEN_7396; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_br = slots_18_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7595 = _T_965 ? issue_slots_18_uop_is_br : _GEN_7397; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_iw_p2_poisoned = slots_18_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7596 = _T_965 ? issue_slots_18_uop_iw_p2_poisoned : _GEN_7398; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_iw_p1_poisoned = slots_18_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7597 = _T_965 ? issue_slots_18_uop_iw_p1_poisoned : _GEN_7399; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_iw_state = slots_18_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7598 = _T_965 ? issue_slots_18_uop_iw_state : _GEN_7400; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_ctrl_op3_sel = slots_18_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7599 = _T_965 ? issue_slots_18_uop_ctrl_op3_sel : _GEN_7401; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_ctrl_is_std = slots_18_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7600 = _T_965 ? issue_slots_18_uop_ctrl_is_std : _GEN_7402; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_ctrl_is_sta = slots_18_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7601 = _T_965 ? issue_slots_18_uop_ctrl_is_sta : _GEN_7403; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_ctrl_is_load = slots_18_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7602 = _T_965 ? issue_slots_18_uop_ctrl_is_load : _GEN_7404; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_18_uop_ctrl_csr_cmd = slots_18_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7603 = _T_965 ? issue_slots_18_uop_ctrl_csr_cmd : _GEN_7405; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_ctrl_fcn_dw = slots_18_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7604 = _T_965 ? issue_slots_18_uop_ctrl_fcn_dw : _GEN_7406; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_ctrl_op_fcn = slots_18_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7605 = _T_965 ? issue_slots_18_uop_ctrl_op_fcn : _GEN_7407; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_18_uop_ctrl_imm_sel = slots_18_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7606 = _T_965 ? issue_slots_18_uop_ctrl_imm_sel : _GEN_7408; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_18_uop_ctrl_op2_sel = slots_18_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7607 = _T_965 ? issue_slots_18_uop_ctrl_op2_sel : _GEN_7409; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_ctrl_op1_sel = slots_18_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7608 = _T_965 ? issue_slots_18_uop_ctrl_op1_sel : _GEN_7410; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_ctrl_br_type = slots_18_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7609 = _T_965 ? issue_slots_18_uop_ctrl_br_type : _GEN_7411; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7610 = _T_965 ? issue_slots_18_uop_fu_code : _GEN_7412; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_18_uop_iq_type = slots_18_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7611 = _T_965 ? issue_slots_18_uop_iq_type : _GEN_7413; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_18_uop_debug_pc = slots_18_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_7612 = _T_965 ? issue_slots_18_uop_debug_pc : _GEN_7414; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_rvc = slots_18_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7613 = _T_965 ? issue_slots_18_uop_is_rvc : _GEN_7415; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_18_uop_debug_inst = slots_18_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7614 = _T_965 ? issue_slots_18_uop_debug_inst : _GEN_7416; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_18_uop_inst = slots_18_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_7615 = _T_965 ? issue_slots_18_uop_inst : _GEN_7417; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_18_uop_uopc = slots_18_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_7616 = _T_965 ? issue_slots_18_uop_uopc : _GEN_7418; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_address_num = slots_18_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7617 = _T_965 ? issue_slots_18_uop_address_num : _GEN_7419; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_rob_inst_idx = slots_18_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7618 = _T_965 ? issue_slots_18_uop_rob_inst_idx : _GEN_7420; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_self_index = slots_18_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7619 = _T_965 ? issue_slots_18_uop_self_index : _GEN_7421; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_18_uop_split_num = slots_18_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_7620 = _T_965 ? issue_slots_18_uop_split_num : _GEN_7422; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_op2_sel = slots_18_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7621 = _T_965 ? issue_slots_18_uop_op2_sel : _GEN_7423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_op1_sel = slots_18_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7622 = _T_965 ? issue_slots_18_uop_op1_sel : _GEN_7424; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_stale_pflag = slots_18_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7623 = _T_965 ? issue_slots_18_uop_stale_pflag : _GEN_7425; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_pflag_busy = slots_18_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7624 = _T_965 ? issue_slots_18_uop_pflag_busy : _GEN_7426; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_pwflag = slots_18_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7625 = _T_965 ? issue_slots_18_uop_pwflag : _GEN_7427; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_18_uop_prflag = slots_18_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_7626 = _T_965 ? issue_slots_18_uop_prflag : _GEN_7428; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_wflag = slots_18_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7627 = _T_965 ? issue_slots_18_uop_wflag : _GEN_7429; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_rflag = slots_18_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7628 = _T_965 ? issue_slots_18_uop_rflag : _GEN_7430; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_18_uop_lrs3_rtype = slots_18_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_7629 = _T_965 ? issue_slots_18_uop_lrs3_rtype : _GEN_7431; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_18_uop_shift = slots_18_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_7630 = _T_965 ? issue_slots_18_uop_shift : _GEN_7432; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_is_unicore = slots_18_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7631 = _T_965 ? issue_slots_18_uop_is_unicore : _GEN_7433; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_switch_off = slots_18_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7632 = _T_965 ? issue_slots_18_uop_switch_off : _GEN_7434; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_18_uop_switch = slots_18_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_7633 = _T_965 ? issue_slots_18_uop_switch : _GEN_7435; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7636 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_debug_tsrc : _GEN_7438
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7637 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_debug_fsrc : _GEN_7439
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7638 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_bp_xcpt_if : _GEN_7440; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7639 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_bp_debug_if : _GEN_7441; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7640 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_xcpt_ma_if : _GEN_7442; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7641 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_xcpt_ae_if : _GEN_7443; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7642 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_xcpt_pf_if : _GEN_7444; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7643 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_fp_single : _GEN_7445; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7644 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_fp_val : _GEN_7446; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7645 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_frs3_en : _GEN_7447; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7646 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_lrs2_rtype : _GEN_7448
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7647 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_lrs1_rtype : _GEN_7449
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7648 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_dst_rtype : _GEN_7450; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7649 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ldst_val : _GEN_7451; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7650 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_lrs3 : _GEN_7452; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7651 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_lrs2 : _GEN_7453; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7652 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_lrs1 : _GEN_7454; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7653 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ldst : _GEN_7455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7654 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ldst_is_rs1 : _GEN_7456; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7655 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_flush_on_commit : _GEN_7457
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7656 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_unique : _GEN_7458; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7657 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_sys_pc2epc : _GEN_7459; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7658 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_uses_stq : _GEN_7460; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7659 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_uses_ldq : _GEN_7461; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7660 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_amo : _GEN_7462; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7661 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_fencei : _GEN_7463; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7662 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_fence : _GEN_7464; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7663 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_mem_signed : _GEN_7465; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7664 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_mem_size : _GEN_7466; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7665 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_mem_cmd : _GEN_7467; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7666 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_bypassable : _GEN_7468; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] _GEN_7667 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_exc_cause : _GEN_7469
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7668 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_exception : _GEN_7470; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7669 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_stale_pdst : _GEN_7471
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7670 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ppred_busy : _GEN_7472; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7671 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_prs3_busy : _GEN_7473; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7672 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_prs2_busy : _GEN_7474; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7673 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_prs1_busy : _GEN_7475; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7674 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ppred : _GEN_7476; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7675 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_prs3 : _GEN_7477; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7676 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_prs2 : _GEN_7478; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7677 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_prs1 : _GEN_7479; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7678 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_pdst : _GEN_7480; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7679 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_rxq_idx : _GEN_7481; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7680 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_stq_idx : _GEN_7482; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7681 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ldq_idx : _GEN_7483; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7682 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_rob_idx : _GEN_7484; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7683 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_csr_addr : _GEN_7485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] _GEN_7684 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_imm_packed :
    _GEN_7486; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7685 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_taken : _GEN_7487; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7686 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_pc_lob : _GEN_7488; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7687 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_edge_inst : _GEN_7489; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] _GEN_7688 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ftq_idx : _GEN_7490; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7689 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_br_tag : _GEN_7491; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] _GEN_7690 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_br_mask : _GEN_7492; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7691 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_sfb : _GEN_7493; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7692 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_jal : _GEN_7494; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7693 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_jalr : _GEN_7495; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7694 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_br : _GEN_7496; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7695 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_iw_p2_poisoned : _GEN_7497; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7696 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_iw_p1_poisoned : _GEN_7498; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7697 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_iw_state : _GEN_7499; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7698 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_op3_sel :
    _GEN_7500; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7699 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_is_std : _GEN_7501; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7700 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_is_sta : _GEN_7502; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7701 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_is_load : _GEN_7503; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7702 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_csr_cmd :
    _GEN_7504; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7703 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_fcn_dw : _GEN_7505; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7704 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_op_fcn :
    _GEN_7506; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7705 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_imm_sel :
    _GEN_7507; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7706 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_op2_sel :
    _GEN_7508; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7707 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_op1_sel :
    _GEN_7509; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7708 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_ctrl_br_type :
    _GEN_7510; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_7709 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_fu_code : _GEN_7511; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7710 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_iq_type : _GEN_7512; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] _GEN_7711 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_debug_pc : _GEN_7513; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7712 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_rvc : _GEN_7514; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7713 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_debug_inst :
    _GEN_7515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] _GEN_7714 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_inst : _GEN_7516; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] _GEN_7715 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_uopc : _GEN_7517; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7716 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_address_num :
    _GEN_7518; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7717 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_rob_inst_idx :
    _GEN_7519; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7718 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_self_index : _GEN_7520
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] _GEN_7719 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_split_num : _GEN_7521; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7720 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_op2_sel : _GEN_7522; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7721 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_op1_sel : _GEN_7523; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7722 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_stale_pflag :
    _GEN_7524; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7723 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_pflag_busy : _GEN_7525; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7724 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_pwflag : _GEN_7526; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] _GEN_7725 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_prflag : _GEN_7527; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7726 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_wflag : _GEN_7528; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7727 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_rflag : _GEN_7529; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] _GEN_7728 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_lrs3_rtype : _GEN_7530
    ; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] _GEN_7729 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_shift : _GEN_7531; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7730 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_is_unicore : _GEN_7532; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7731 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_switch_off : _GEN_7533; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  _GEN_7732 = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 ? issue_slots_18_uop_switch : _GEN_7534; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_19_uop_debug_tsrc = slots_19_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_debug_fsrc = slots_19_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_bp_xcpt_if = slots_19_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_bp_debug_if = slots_19_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_xcpt_ma_if = slots_19_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_xcpt_ae_if = slots_19_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_xcpt_pf_if = slots_19_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_fp_single = slots_19_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_fp_val = slots_19_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_frs3_en = slots_19_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_lrs2_rtype = slots_19_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_lrs1_rtype = slots_19_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_dst_rtype = slots_19_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_ldst_val = slots_19_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_lrs3 = slots_19_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_lrs2 = slots_19_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_lrs1 = slots_19_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_ldst = slots_19_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_ldst_is_rs1 = slots_19_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_flush_on_commit = slots_19_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_unique = slots_19_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_sys_pc2epc = slots_19_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_uses_stq = slots_19_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_uses_ldq = slots_19_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_amo = slots_19_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_fencei = slots_19_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_fence = slots_19_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_mem_signed = slots_19_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_mem_size = slots_19_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_uop_mem_cmd = slots_19_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_bypassable = slots_19_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_19_uop_exc_cause = slots_19_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_exception = slots_19_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_uop_stale_pdst = slots_19_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_ppred_busy = slots_19_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_prs3_busy = slots_19_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_prs2_busy = slots_19_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_prs1_busy = slots_19_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_uop_ppred = slots_19_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_uop_prs3 = slots_19_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_uop_prs2 = slots_19_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_uop_prs1 = slots_19_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_uop_pdst = slots_19_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_rxq_idx = slots_19_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_uop_stq_idx = slots_19_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_uop_ldq_idx = slots_19_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_rob_idx = slots_19_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_19_uop_csr_addr = slots_19_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_19_uop_imm_packed = slots_19_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_taken = slots_19_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_pc_lob = slots_19_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_edge_inst = slots_19_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_19_uop_ftq_idx = slots_19_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_br_tag = slots_19_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_19_uop_br_mask = slots_19_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_sfb = slots_19_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_jal = slots_19_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_jalr = slots_19_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_br = slots_19_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_iw_p2_poisoned = slots_19_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_iw_p1_poisoned = slots_19_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_iw_state = slots_19_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_ctrl_op3_sel = slots_19_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_ctrl_is_std = slots_19_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_ctrl_is_sta = slots_19_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_ctrl_is_load = slots_19_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_uop_ctrl_csr_cmd = slots_19_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_ctrl_fcn_dw = slots_19_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_ctrl_op_fcn = slots_19_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_uop_ctrl_imm_sel = slots_19_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_uop_ctrl_op2_sel = slots_19_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_ctrl_op1_sel = slots_19_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_ctrl_br_type = slots_19_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_uop_iq_type = slots_19_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_19_uop_debug_pc = slots_19_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_rvc = slots_19_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_19_uop_debug_inst = slots_19_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_19_uop_inst = slots_19_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_19_uop_uopc = slots_19_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_address_num = slots_19_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_rob_inst_idx = slots_19_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_self_index = slots_19_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_19_uop_split_num = slots_19_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_op2_sel = slots_19_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_op1_sel = slots_19_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_stale_pflag = slots_19_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_pflag_busy = slots_19_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_pwflag = slots_19_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_19_uop_prflag = slots_19_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_wflag = slots_19_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_rflag = slots_19_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_19_uop_lrs3_rtype = slots_19_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_19_uop_shift = slots_19_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_is_unicore = slots_19_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_switch_off = slots_19_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_19_uop_switch = slots_19_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  IssueSlot_16 slots_0 ( // @[issue-unit.scala 157:73]
    .clock(slots_0_clock),
    .reset(slots_0_reset),
    .io_valid(slots_0_io_valid),
    .io_will_be_valid(slots_0_io_will_be_valid),
    .io_request(slots_0_io_request),
    .io_request_hp(slots_0_io_request_hp),
    .io_grant(slots_0_io_grant),
    .io_brupdate_b1_resolve_mask(slots_0_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_0_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_0_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_0_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_0_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_0_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_0_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_0_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_0_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_0_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_0_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_0_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_0_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_0_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_0_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_0_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_0_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_0_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_0_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_0_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_0_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_0_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_0_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_0_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_0_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_0_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_0_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_0_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_0_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_0_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_0_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_0_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_0_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_0_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_0_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_0_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_0_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_0_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_0_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_0_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_0_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_0_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_0_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_0_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_0_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_0_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_0_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_0_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_0_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_0_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_0_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_0_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_0_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_0_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_0_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_0_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_0_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_0_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_0_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_0_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_0_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_0_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_0_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_0_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_0_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_0_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_0_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_0_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_0_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_0_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_0_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_0_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_0_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_0_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_0_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_0_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_0_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_0_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_0_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_0_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_0_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_0_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_0_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_0_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_0_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_0_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_0_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_0_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_0_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_0_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_0_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_0_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_0_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_0_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_0_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_0_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_0_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_0_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_0_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_0_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_0_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_0_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_0_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_0_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_0_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_0_io_brupdate_b2_target_offset),
    .io_kill(slots_0_io_kill),
    .io_clear(slots_0_io_clear),
    .io_ldspec_miss(slots_0_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_0_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_0_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_0_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_0_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_0_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_0_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_0_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_0_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_0_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_0_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_0_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_0_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_0_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_0_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_0_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_0_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_0_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_0_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_0_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_0_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_0_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_0_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_0_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_0_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_0_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_0_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_0_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_0_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_0_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_0_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_0_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_0_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_0_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_0_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_0_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_0_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_0_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_0_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_0_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_0_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_0_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_0_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_0_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_0_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_0_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_0_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_0_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_0_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_0_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_0_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_0_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_0_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_0_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_0_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_0_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_0_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_0_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_0_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_0_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_0_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_0_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_0_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_0_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_0_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_0_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_0_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_0_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_0_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_0_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_0_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_0_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_0_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_0_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_0_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_0_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_0_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_0_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_0_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_0_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_0_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_0_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_0_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_0_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_0_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_0_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_0_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_0_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_0_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_0_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_0_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_0_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_0_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_0_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_0_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_0_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_0_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_0_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_0_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_0_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_0_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_0_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_0_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_0_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_0_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_0_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_0_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_0_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_0_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_0_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_0_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_0_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_0_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_0_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_0_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_0_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_0_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_0_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_0_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_0_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_0_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_0_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_0_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_0_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_0_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_0_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_0_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_0_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_0_io_out_uop_switch),
    .io_out_uop_switch_off(slots_0_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_0_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_0_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_0_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_0_io_out_uop_rflag),
    .io_out_uop_wflag(slots_0_io_out_uop_wflag),
    .io_out_uop_prflag(slots_0_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_0_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_0_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_0_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_0_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_0_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_0_io_out_uop_split_num),
    .io_out_uop_self_index(slots_0_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_0_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_0_io_out_uop_address_num),
    .io_out_uop_uopc(slots_0_io_out_uop_uopc),
    .io_out_uop_inst(slots_0_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_0_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_0_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_0_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_0_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_0_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_0_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_0_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_0_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_0_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_0_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_0_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_0_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_0_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_0_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_0_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_0_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_0_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_0_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_0_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_0_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_0_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_0_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_0_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_0_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_0_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_0_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_0_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_0_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_0_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_0_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_0_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_0_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_0_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_0_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_0_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_0_io_out_uop_pdst),
    .io_out_uop_prs1(slots_0_io_out_uop_prs1),
    .io_out_uop_prs2(slots_0_io_out_uop_prs2),
    .io_out_uop_prs3(slots_0_io_out_uop_prs3),
    .io_out_uop_ppred(slots_0_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_0_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_0_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_0_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_0_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_0_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_0_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_0_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_0_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_0_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_0_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_0_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_0_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_0_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_0_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_0_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_0_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_0_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_0_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_0_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_0_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_0_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_0_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_0_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_0_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_0_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_0_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_0_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_0_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_0_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_0_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_0_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_0_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_0_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_0_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_0_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_0_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_0_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_0_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_0_io_uop_switch),
    .io_uop_switch_off(slots_0_io_uop_switch_off),
    .io_uop_is_unicore(slots_0_io_uop_is_unicore),
    .io_uop_shift(slots_0_io_uop_shift),
    .io_uop_lrs3_rtype(slots_0_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_0_io_uop_rflag),
    .io_uop_wflag(slots_0_io_uop_wflag),
    .io_uop_prflag(slots_0_io_uop_prflag),
    .io_uop_pwflag(slots_0_io_uop_pwflag),
    .io_uop_pflag_busy(slots_0_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_0_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_0_io_uop_op1_sel),
    .io_uop_op2_sel(slots_0_io_uop_op2_sel),
    .io_uop_split_num(slots_0_io_uop_split_num),
    .io_uop_self_index(slots_0_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_0_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_0_io_uop_address_num),
    .io_uop_uopc(slots_0_io_uop_uopc),
    .io_uop_inst(slots_0_io_uop_inst),
    .io_uop_debug_inst(slots_0_io_uop_debug_inst),
    .io_uop_is_rvc(slots_0_io_uop_is_rvc),
    .io_uop_debug_pc(slots_0_io_uop_debug_pc),
    .io_uop_iq_type(slots_0_io_uop_iq_type),
    .io_uop_fu_code(slots_0_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_0_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_0_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_0_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_0_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_0_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_0_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_0_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_0_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_0_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_0_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_0_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_0_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_0_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_0_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_0_io_uop_is_br),
    .io_uop_is_jalr(slots_0_io_uop_is_jalr),
    .io_uop_is_jal(slots_0_io_uop_is_jal),
    .io_uop_is_sfb(slots_0_io_uop_is_sfb),
    .io_uop_br_mask(slots_0_io_uop_br_mask),
    .io_uop_br_tag(slots_0_io_uop_br_tag),
    .io_uop_ftq_idx(slots_0_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_0_io_uop_edge_inst),
    .io_uop_pc_lob(slots_0_io_uop_pc_lob),
    .io_uop_taken(slots_0_io_uop_taken),
    .io_uop_imm_packed(slots_0_io_uop_imm_packed),
    .io_uop_csr_addr(slots_0_io_uop_csr_addr),
    .io_uop_rob_idx(slots_0_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_0_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_0_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_0_io_uop_rxq_idx),
    .io_uop_pdst(slots_0_io_uop_pdst),
    .io_uop_prs1(slots_0_io_uop_prs1),
    .io_uop_prs2(slots_0_io_uop_prs2),
    .io_uop_prs3(slots_0_io_uop_prs3),
    .io_uop_ppred(slots_0_io_uop_ppred),
    .io_uop_prs1_busy(slots_0_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_0_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_0_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_0_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_0_io_uop_stale_pdst),
    .io_uop_exception(slots_0_io_uop_exception),
    .io_uop_exc_cause(slots_0_io_uop_exc_cause),
    .io_uop_bypassable(slots_0_io_uop_bypassable),
    .io_uop_mem_cmd(slots_0_io_uop_mem_cmd),
    .io_uop_mem_size(slots_0_io_uop_mem_size),
    .io_uop_mem_signed(slots_0_io_uop_mem_signed),
    .io_uop_is_fence(slots_0_io_uop_is_fence),
    .io_uop_is_fencei(slots_0_io_uop_is_fencei),
    .io_uop_is_amo(slots_0_io_uop_is_amo),
    .io_uop_uses_ldq(slots_0_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_0_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_0_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_0_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_0_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_0_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_0_io_uop_ldst),
    .io_uop_lrs1(slots_0_io_uop_lrs1),
    .io_uop_lrs2(slots_0_io_uop_lrs2),
    .io_uop_lrs3(slots_0_io_uop_lrs3),
    .io_uop_ldst_val(slots_0_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_0_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_0_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_0_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_0_io_uop_frs3_en),
    .io_uop_fp_val(slots_0_io_uop_fp_val),
    .io_uop_fp_single(slots_0_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_0_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_0_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_0_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_0_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_0_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_0_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_0_io_uop_debug_tsrc),
    .io_debug_p1(slots_0_io_debug_p1),
    .io_debug_p2(slots_0_io_debug_p2),
    .io_debug_p3(slots_0_io_debug_p3),
    .io_debug_ppred(slots_0_io_debug_ppred),
    .io_debug_state(slots_0_io_debug_state)
  );
  IssueSlot_16 slots_1 ( // @[issue-unit.scala 157:73]
    .clock(slots_1_clock),
    .reset(slots_1_reset),
    .io_valid(slots_1_io_valid),
    .io_will_be_valid(slots_1_io_will_be_valid),
    .io_request(slots_1_io_request),
    .io_request_hp(slots_1_io_request_hp),
    .io_grant(slots_1_io_grant),
    .io_brupdate_b1_resolve_mask(slots_1_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_1_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_1_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_1_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_1_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_1_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_1_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_1_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_1_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_1_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_1_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_1_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_1_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_1_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_1_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_1_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_1_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_1_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_1_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_1_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_1_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_1_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_1_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_1_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_1_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_1_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_1_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_1_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_1_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_1_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_1_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_1_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_1_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_1_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_1_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_1_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_1_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_1_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_1_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_1_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_1_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_1_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_1_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_1_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_1_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_1_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_1_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_1_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_1_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_1_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_1_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_1_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_1_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_1_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_1_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_1_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_1_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_1_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_1_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_1_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_1_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_1_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_1_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_1_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_1_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_1_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_1_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_1_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_1_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_1_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_1_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_1_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_1_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_1_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_1_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_1_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_1_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_1_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_1_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_1_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_1_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_1_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_1_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_1_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_1_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_1_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_1_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_1_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_1_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_1_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_1_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_1_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_1_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_1_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_1_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_1_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_1_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_1_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_1_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_1_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_1_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_1_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_1_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_1_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_1_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_1_io_brupdate_b2_target_offset),
    .io_kill(slots_1_io_kill),
    .io_clear(slots_1_io_clear),
    .io_ldspec_miss(slots_1_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_1_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_1_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_1_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_1_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_1_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_1_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_1_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_1_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_1_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_1_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_1_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_1_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_1_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_1_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_1_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_1_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_1_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_1_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_1_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_1_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_1_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_1_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_1_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_1_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_1_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_1_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_1_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_1_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_1_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_1_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_1_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_1_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_1_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_1_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_1_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_1_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_1_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_1_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_1_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_1_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_1_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_1_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_1_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_1_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_1_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_1_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_1_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_1_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_1_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_1_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_1_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_1_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_1_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_1_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_1_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_1_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_1_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_1_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_1_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_1_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_1_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_1_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_1_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_1_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_1_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_1_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_1_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_1_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_1_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_1_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_1_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_1_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_1_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_1_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_1_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_1_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_1_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_1_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_1_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_1_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_1_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_1_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_1_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_1_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_1_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_1_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_1_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_1_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_1_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_1_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_1_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_1_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_1_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_1_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_1_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_1_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_1_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_1_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_1_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_1_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_1_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_1_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_1_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_1_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_1_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_1_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_1_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_1_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_1_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_1_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_1_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_1_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_1_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_1_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_1_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_1_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_1_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_1_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_1_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_1_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_1_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_1_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_1_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_1_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_1_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_1_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_1_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_1_io_out_uop_switch),
    .io_out_uop_switch_off(slots_1_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_1_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_1_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_1_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_1_io_out_uop_rflag),
    .io_out_uop_wflag(slots_1_io_out_uop_wflag),
    .io_out_uop_prflag(slots_1_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_1_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_1_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_1_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_1_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_1_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_1_io_out_uop_split_num),
    .io_out_uop_self_index(slots_1_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_1_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_1_io_out_uop_address_num),
    .io_out_uop_uopc(slots_1_io_out_uop_uopc),
    .io_out_uop_inst(slots_1_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_1_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_1_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_1_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_1_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_1_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_1_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_1_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_1_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_1_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_1_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_1_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_1_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_1_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_1_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_1_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_1_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_1_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_1_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_1_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_1_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_1_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_1_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_1_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_1_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_1_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_1_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_1_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_1_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_1_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_1_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_1_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_1_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_1_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_1_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_1_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_1_io_out_uop_pdst),
    .io_out_uop_prs1(slots_1_io_out_uop_prs1),
    .io_out_uop_prs2(slots_1_io_out_uop_prs2),
    .io_out_uop_prs3(slots_1_io_out_uop_prs3),
    .io_out_uop_ppred(slots_1_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_1_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_1_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_1_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_1_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_1_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_1_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_1_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_1_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_1_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_1_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_1_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_1_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_1_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_1_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_1_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_1_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_1_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_1_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_1_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_1_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_1_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_1_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_1_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_1_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_1_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_1_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_1_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_1_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_1_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_1_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_1_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_1_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_1_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_1_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_1_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_1_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_1_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_1_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_1_io_uop_switch),
    .io_uop_switch_off(slots_1_io_uop_switch_off),
    .io_uop_is_unicore(slots_1_io_uop_is_unicore),
    .io_uop_shift(slots_1_io_uop_shift),
    .io_uop_lrs3_rtype(slots_1_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_1_io_uop_rflag),
    .io_uop_wflag(slots_1_io_uop_wflag),
    .io_uop_prflag(slots_1_io_uop_prflag),
    .io_uop_pwflag(slots_1_io_uop_pwflag),
    .io_uop_pflag_busy(slots_1_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_1_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_1_io_uop_op1_sel),
    .io_uop_op2_sel(slots_1_io_uop_op2_sel),
    .io_uop_split_num(slots_1_io_uop_split_num),
    .io_uop_self_index(slots_1_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_1_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_1_io_uop_address_num),
    .io_uop_uopc(slots_1_io_uop_uopc),
    .io_uop_inst(slots_1_io_uop_inst),
    .io_uop_debug_inst(slots_1_io_uop_debug_inst),
    .io_uop_is_rvc(slots_1_io_uop_is_rvc),
    .io_uop_debug_pc(slots_1_io_uop_debug_pc),
    .io_uop_iq_type(slots_1_io_uop_iq_type),
    .io_uop_fu_code(slots_1_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_1_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_1_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_1_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_1_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_1_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_1_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_1_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_1_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_1_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_1_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_1_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_1_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_1_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_1_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_1_io_uop_is_br),
    .io_uop_is_jalr(slots_1_io_uop_is_jalr),
    .io_uop_is_jal(slots_1_io_uop_is_jal),
    .io_uop_is_sfb(slots_1_io_uop_is_sfb),
    .io_uop_br_mask(slots_1_io_uop_br_mask),
    .io_uop_br_tag(slots_1_io_uop_br_tag),
    .io_uop_ftq_idx(slots_1_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_1_io_uop_edge_inst),
    .io_uop_pc_lob(slots_1_io_uop_pc_lob),
    .io_uop_taken(slots_1_io_uop_taken),
    .io_uop_imm_packed(slots_1_io_uop_imm_packed),
    .io_uop_csr_addr(slots_1_io_uop_csr_addr),
    .io_uop_rob_idx(slots_1_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_1_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_1_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_1_io_uop_rxq_idx),
    .io_uop_pdst(slots_1_io_uop_pdst),
    .io_uop_prs1(slots_1_io_uop_prs1),
    .io_uop_prs2(slots_1_io_uop_prs2),
    .io_uop_prs3(slots_1_io_uop_prs3),
    .io_uop_ppred(slots_1_io_uop_ppred),
    .io_uop_prs1_busy(slots_1_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_1_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_1_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_1_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_1_io_uop_stale_pdst),
    .io_uop_exception(slots_1_io_uop_exception),
    .io_uop_exc_cause(slots_1_io_uop_exc_cause),
    .io_uop_bypassable(slots_1_io_uop_bypassable),
    .io_uop_mem_cmd(slots_1_io_uop_mem_cmd),
    .io_uop_mem_size(slots_1_io_uop_mem_size),
    .io_uop_mem_signed(slots_1_io_uop_mem_signed),
    .io_uop_is_fence(slots_1_io_uop_is_fence),
    .io_uop_is_fencei(slots_1_io_uop_is_fencei),
    .io_uop_is_amo(slots_1_io_uop_is_amo),
    .io_uop_uses_ldq(slots_1_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_1_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_1_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_1_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_1_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_1_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_1_io_uop_ldst),
    .io_uop_lrs1(slots_1_io_uop_lrs1),
    .io_uop_lrs2(slots_1_io_uop_lrs2),
    .io_uop_lrs3(slots_1_io_uop_lrs3),
    .io_uop_ldst_val(slots_1_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_1_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_1_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_1_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_1_io_uop_frs3_en),
    .io_uop_fp_val(slots_1_io_uop_fp_val),
    .io_uop_fp_single(slots_1_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_1_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_1_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_1_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_1_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_1_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_1_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_1_io_uop_debug_tsrc),
    .io_debug_p1(slots_1_io_debug_p1),
    .io_debug_p2(slots_1_io_debug_p2),
    .io_debug_p3(slots_1_io_debug_p3),
    .io_debug_ppred(slots_1_io_debug_ppred),
    .io_debug_state(slots_1_io_debug_state)
  );
  IssueSlot_16 slots_2 ( // @[issue-unit.scala 157:73]
    .clock(slots_2_clock),
    .reset(slots_2_reset),
    .io_valid(slots_2_io_valid),
    .io_will_be_valid(slots_2_io_will_be_valid),
    .io_request(slots_2_io_request),
    .io_request_hp(slots_2_io_request_hp),
    .io_grant(slots_2_io_grant),
    .io_brupdate_b1_resolve_mask(slots_2_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_2_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_2_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_2_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_2_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_2_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_2_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_2_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_2_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_2_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_2_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_2_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_2_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_2_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_2_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_2_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_2_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_2_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_2_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_2_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_2_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_2_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_2_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_2_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_2_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_2_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_2_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_2_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_2_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_2_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_2_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_2_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_2_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_2_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_2_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_2_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_2_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_2_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_2_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_2_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_2_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_2_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_2_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_2_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_2_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_2_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_2_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_2_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_2_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_2_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_2_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_2_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_2_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_2_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_2_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_2_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_2_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_2_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_2_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_2_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_2_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_2_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_2_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_2_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_2_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_2_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_2_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_2_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_2_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_2_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_2_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_2_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_2_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_2_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_2_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_2_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_2_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_2_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_2_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_2_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_2_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_2_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_2_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_2_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_2_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_2_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_2_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_2_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_2_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_2_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_2_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_2_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_2_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_2_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_2_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_2_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_2_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_2_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_2_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_2_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_2_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_2_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_2_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_2_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_2_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_2_io_brupdate_b2_target_offset),
    .io_kill(slots_2_io_kill),
    .io_clear(slots_2_io_clear),
    .io_ldspec_miss(slots_2_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_2_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_2_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_2_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_2_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_2_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_2_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_2_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_2_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_2_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_2_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_2_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_2_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_2_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_2_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_2_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_2_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_2_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_2_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_2_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_2_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_2_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_2_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_2_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_2_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_2_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_2_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_2_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_2_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_2_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_2_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_2_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_2_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_2_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_2_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_2_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_2_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_2_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_2_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_2_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_2_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_2_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_2_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_2_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_2_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_2_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_2_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_2_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_2_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_2_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_2_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_2_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_2_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_2_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_2_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_2_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_2_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_2_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_2_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_2_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_2_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_2_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_2_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_2_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_2_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_2_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_2_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_2_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_2_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_2_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_2_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_2_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_2_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_2_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_2_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_2_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_2_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_2_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_2_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_2_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_2_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_2_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_2_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_2_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_2_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_2_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_2_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_2_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_2_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_2_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_2_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_2_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_2_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_2_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_2_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_2_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_2_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_2_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_2_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_2_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_2_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_2_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_2_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_2_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_2_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_2_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_2_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_2_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_2_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_2_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_2_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_2_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_2_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_2_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_2_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_2_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_2_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_2_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_2_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_2_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_2_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_2_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_2_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_2_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_2_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_2_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_2_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_2_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_2_io_out_uop_switch),
    .io_out_uop_switch_off(slots_2_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_2_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_2_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_2_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_2_io_out_uop_rflag),
    .io_out_uop_wflag(slots_2_io_out_uop_wflag),
    .io_out_uop_prflag(slots_2_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_2_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_2_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_2_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_2_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_2_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_2_io_out_uop_split_num),
    .io_out_uop_self_index(slots_2_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_2_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_2_io_out_uop_address_num),
    .io_out_uop_uopc(slots_2_io_out_uop_uopc),
    .io_out_uop_inst(slots_2_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_2_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_2_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_2_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_2_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_2_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_2_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_2_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_2_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_2_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_2_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_2_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_2_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_2_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_2_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_2_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_2_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_2_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_2_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_2_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_2_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_2_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_2_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_2_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_2_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_2_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_2_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_2_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_2_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_2_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_2_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_2_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_2_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_2_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_2_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_2_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_2_io_out_uop_pdst),
    .io_out_uop_prs1(slots_2_io_out_uop_prs1),
    .io_out_uop_prs2(slots_2_io_out_uop_prs2),
    .io_out_uop_prs3(slots_2_io_out_uop_prs3),
    .io_out_uop_ppred(slots_2_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_2_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_2_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_2_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_2_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_2_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_2_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_2_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_2_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_2_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_2_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_2_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_2_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_2_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_2_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_2_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_2_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_2_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_2_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_2_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_2_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_2_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_2_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_2_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_2_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_2_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_2_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_2_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_2_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_2_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_2_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_2_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_2_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_2_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_2_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_2_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_2_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_2_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_2_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_2_io_uop_switch),
    .io_uop_switch_off(slots_2_io_uop_switch_off),
    .io_uop_is_unicore(slots_2_io_uop_is_unicore),
    .io_uop_shift(slots_2_io_uop_shift),
    .io_uop_lrs3_rtype(slots_2_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_2_io_uop_rflag),
    .io_uop_wflag(slots_2_io_uop_wflag),
    .io_uop_prflag(slots_2_io_uop_prflag),
    .io_uop_pwflag(slots_2_io_uop_pwflag),
    .io_uop_pflag_busy(slots_2_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_2_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_2_io_uop_op1_sel),
    .io_uop_op2_sel(slots_2_io_uop_op2_sel),
    .io_uop_split_num(slots_2_io_uop_split_num),
    .io_uop_self_index(slots_2_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_2_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_2_io_uop_address_num),
    .io_uop_uopc(slots_2_io_uop_uopc),
    .io_uop_inst(slots_2_io_uop_inst),
    .io_uop_debug_inst(slots_2_io_uop_debug_inst),
    .io_uop_is_rvc(slots_2_io_uop_is_rvc),
    .io_uop_debug_pc(slots_2_io_uop_debug_pc),
    .io_uop_iq_type(slots_2_io_uop_iq_type),
    .io_uop_fu_code(slots_2_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_2_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_2_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_2_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_2_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_2_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_2_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_2_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_2_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_2_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_2_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_2_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_2_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_2_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_2_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_2_io_uop_is_br),
    .io_uop_is_jalr(slots_2_io_uop_is_jalr),
    .io_uop_is_jal(slots_2_io_uop_is_jal),
    .io_uop_is_sfb(slots_2_io_uop_is_sfb),
    .io_uop_br_mask(slots_2_io_uop_br_mask),
    .io_uop_br_tag(slots_2_io_uop_br_tag),
    .io_uop_ftq_idx(slots_2_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_2_io_uop_edge_inst),
    .io_uop_pc_lob(slots_2_io_uop_pc_lob),
    .io_uop_taken(slots_2_io_uop_taken),
    .io_uop_imm_packed(slots_2_io_uop_imm_packed),
    .io_uop_csr_addr(slots_2_io_uop_csr_addr),
    .io_uop_rob_idx(slots_2_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_2_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_2_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_2_io_uop_rxq_idx),
    .io_uop_pdst(slots_2_io_uop_pdst),
    .io_uop_prs1(slots_2_io_uop_prs1),
    .io_uop_prs2(slots_2_io_uop_prs2),
    .io_uop_prs3(slots_2_io_uop_prs3),
    .io_uop_ppred(slots_2_io_uop_ppred),
    .io_uop_prs1_busy(slots_2_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_2_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_2_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_2_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_2_io_uop_stale_pdst),
    .io_uop_exception(slots_2_io_uop_exception),
    .io_uop_exc_cause(slots_2_io_uop_exc_cause),
    .io_uop_bypassable(slots_2_io_uop_bypassable),
    .io_uop_mem_cmd(slots_2_io_uop_mem_cmd),
    .io_uop_mem_size(slots_2_io_uop_mem_size),
    .io_uop_mem_signed(slots_2_io_uop_mem_signed),
    .io_uop_is_fence(slots_2_io_uop_is_fence),
    .io_uop_is_fencei(slots_2_io_uop_is_fencei),
    .io_uop_is_amo(slots_2_io_uop_is_amo),
    .io_uop_uses_ldq(slots_2_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_2_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_2_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_2_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_2_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_2_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_2_io_uop_ldst),
    .io_uop_lrs1(slots_2_io_uop_lrs1),
    .io_uop_lrs2(slots_2_io_uop_lrs2),
    .io_uop_lrs3(slots_2_io_uop_lrs3),
    .io_uop_ldst_val(slots_2_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_2_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_2_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_2_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_2_io_uop_frs3_en),
    .io_uop_fp_val(slots_2_io_uop_fp_val),
    .io_uop_fp_single(slots_2_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_2_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_2_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_2_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_2_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_2_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_2_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_2_io_uop_debug_tsrc),
    .io_debug_p1(slots_2_io_debug_p1),
    .io_debug_p2(slots_2_io_debug_p2),
    .io_debug_p3(slots_2_io_debug_p3),
    .io_debug_ppred(slots_2_io_debug_ppred),
    .io_debug_state(slots_2_io_debug_state)
  );
  IssueSlot_16 slots_3 ( // @[issue-unit.scala 157:73]
    .clock(slots_3_clock),
    .reset(slots_3_reset),
    .io_valid(slots_3_io_valid),
    .io_will_be_valid(slots_3_io_will_be_valid),
    .io_request(slots_3_io_request),
    .io_request_hp(slots_3_io_request_hp),
    .io_grant(slots_3_io_grant),
    .io_brupdate_b1_resolve_mask(slots_3_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_3_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_3_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_3_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_3_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_3_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_3_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_3_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_3_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_3_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_3_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_3_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_3_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_3_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_3_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_3_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_3_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_3_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_3_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_3_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_3_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_3_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_3_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_3_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_3_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_3_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_3_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_3_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_3_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_3_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_3_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_3_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_3_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_3_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_3_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_3_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_3_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_3_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_3_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_3_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_3_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_3_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_3_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_3_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_3_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_3_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_3_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_3_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_3_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_3_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_3_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_3_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_3_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_3_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_3_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_3_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_3_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_3_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_3_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_3_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_3_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_3_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_3_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_3_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_3_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_3_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_3_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_3_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_3_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_3_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_3_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_3_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_3_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_3_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_3_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_3_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_3_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_3_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_3_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_3_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_3_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_3_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_3_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_3_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_3_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_3_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_3_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_3_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_3_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_3_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_3_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_3_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_3_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_3_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_3_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_3_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_3_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_3_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_3_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_3_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_3_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_3_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_3_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_3_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_3_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_3_io_brupdate_b2_target_offset),
    .io_kill(slots_3_io_kill),
    .io_clear(slots_3_io_clear),
    .io_ldspec_miss(slots_3_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_3_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_3_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_3_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_3_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_3_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_3_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_3_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_3_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_3_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_3_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_3_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_3_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_3_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_3_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_3_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_3_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_3_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_3_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_3_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_3_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_3_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_3_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_3_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_3_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_3_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_3_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_3_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_3_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_3_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_3_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_3_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_3_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_3_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_3_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_3_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_3_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_3_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_3_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_3_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_3_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_3_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_3_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_3_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_3_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_3_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_3_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_3_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_3_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_3_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_3_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_3_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_3_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_3_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_3_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_3_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_3_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_3_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_3_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_3_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_3_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_3_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_3_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_3_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_3_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_3_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_3_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_3_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_3_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_3_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_3_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_3_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_3_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_3_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_3_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_3_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_3_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_3_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_3_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_3_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_3_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_3_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_3_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_3_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_3_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_3_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_3_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_3_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_3_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_3_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_3_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_3_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_3_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_3_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_3_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_3_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_3_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_3_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_3_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_3_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_3_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_3_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_3_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_3_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_3_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_3_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_3_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_3_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_3_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_3_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_3_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_3_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_3_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_3_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_3_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_3_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_3_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_3_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_3_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_3_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_3_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_3_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_3_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_3_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_3_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_3_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_3_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_3_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_3_io_out_uop_switch),
    .io_out_uop_switch_off(slots_3_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_3_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_3_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_3_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_3_io_out_uop_rflag),
    .io_out_uop_wflag(slots_3_io_out_uop_wflag),
    .io_out_uop_prflag(slots_3_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_3_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_3_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_3_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_3_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_3_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_3_io_out_uop_split_num),
    .io_out_uop_self_index(slots_3_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_3_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_3_io_out_uop_address_num),
    .io_out_uop_uopc(slots_3_io_out_uop_uopc),
    .io_out_uop_inst(slots_3_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_3_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_3_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_3_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_3_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_3_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_3_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_3_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_3_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_3_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_3_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_3_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_3_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_3_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_3_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_3_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_3_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_3_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_3_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_3_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_3_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_3_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_3_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_3_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_3_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_3_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_3_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_3_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_3_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_3_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_3_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_3_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_3_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_3_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_3_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_3_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_3_io_out_uop_pdst),
    .io_out_uop_prs1(slots_3_io_out_uop_prs1),
    .io_out_uop_prs2(slots_3_io_out_uop_prs2),
    .io_out_uop_prs3(slots_3_io_out_uop_prs3),
    .io_out_uop_ppred(slots_3_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_3_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_3_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_3_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_3_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_3_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_3_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_3_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_3_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_3_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_3_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_3_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_3_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_3_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_3_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_3_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_3_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_3_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_3_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_3_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_3_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_3_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_3_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_3_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_3_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_3_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_3_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_3_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_3_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_3_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_3_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_3_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_3_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_3_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_3_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_3_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_3_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_3_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_3_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_3_io_uop_switch),
    .io_uop_switch_off(slots_3_io_uop_switch_off),
    .io_uop_is_unicore(slots_3_io_uop_is_unicore),
    .io_uop_shift(slots_3_io_uop_shift),
    .io_uop_lrs3_rtype(slots_3_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_3_io_uop_rflag),
    .io_uop_wflag(slots_3_io_uop_wflag),
    .io_uop_prflag(slots_3_io_uop_prflag),
    .io_uop_pwflag(slots_3_io_uop_pwflag),
    .io_uop_pflag_busy(slots_3_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_3_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_3_io_uop_op1_sel),
    .io_uop_op2_sel(slots_3_io_uop_op2_sel),
    .io_uop_split_num(slots_3_io_uop_split_num),
    .io_uop_self_index(slots_3_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_3_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_3_io_uop_address_num),
    .io_uop_uopc(slots_3_io_uop_uopc),
    .io_uop_inst(slots_3_io_uop_inst),
    .io_uop_debug_inst(slots_3_io_uop_debug_inst),
    .io_uop_is_rvc(slots_3_io_uop_is_rvc),
    .io_uop_debug_pc(slots_3_io_uop_debug_pc),
    .io_uop_iq_type(slots_3_io_uop_iq_type),
    .io_uop_fu_code(slots_3_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_3_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_3_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_3_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_3_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_3_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_3_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_3_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_3_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_3_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_3_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_3_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_3_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_3_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_3_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_3_io_uop_is_br),
    .io_uop_is_jalr(slots_3_io_uop_is_jalr),
    .io_uop_is_jal(slots_3_io_uop_is_jal),
    .io_uop_is_sfb(slots_3_io_uop_is_sfb),
    .io_uop_br_mask(slots_3_io_uop_br_mask),
    .io_uop_br_tag(slots_3_io_uop_br_tag),
    .io_uop_ftq_idx(slots_3_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_3_io_uop_edge_inst),
    .io_uop_pc_lob(slots_3_io_uop_pc_lob),
    .io_uop_taken(slots_3_io_uop_taken),
    .io_uop_imm_packed(slots_3_io_uop_imm_packed),
    .io_uop_csr_addr(slots_3_io_uop_csr_addr),
    .io_uop_rob_idx(slots_3_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_3_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_3_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_3_io_uop_rxq_idx),
    .io_uop_pdst(slots_3_io_uop_pdst),
    .io_uop_prs1(slots_3_io_uop_prs1),
    .io_uop_prs2(slots_3_io_uop_prs2),
    .io_uop_prs3(slots_3_io_uop_prs3),
    .io_uop_ppred(slots_3_io_uop_ppred),
    .io_uop_prs1_busy(slots_3_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_3_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_3_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_3_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_3_io_uop_stale_pdst),
    .io_uop_exception(slots_3_io_uop_exception),
    .io_uop_exc_cause(slots_3_io_uop_exc_cause),
    .io_uop_bypassable(slots_3_io_uop_bypassable),
    .io_uop_mem_cmd(slots_3_io_uop_mem_cmd),
    .io_uop_mem_size(slots_3_io_uop_mem_size),
    .io_uop_mem_signed(slots_3_io_uop_mem_signed),
    .io_uop_is_fence(slots_3_io_uop_is_fence),
    .io_uop_is_fencei(slots_3_io_uop_is_fencei),
    .io_uop_is_amo(slots_3_io_uop_is_amo),
    .io_uop_uses_ldq(slots_3_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_3_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_3_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_3_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_3_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_3_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_3_io_uop_ldst),
    .io_uop_lrs1(slots_3_io_uop_lrs1),
    .io_uop_lrs2(slots_3_io_uop_lrs2),
    .io_uop_lrs3(slots_3_io_uop_lrs3),
    .io_uop_ldst_val(slots_3_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_3_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_3_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_3_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_3_io_uop_frs3_en),
    .io_uop_fp_val(slots_3_io_uop_fp_val),
    .io_uop_fp_single(slots_3_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_3_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_3_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_3_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_3_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_3_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_3_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_3_io_uop_debug_tsrc),
    .io_debug_p1(slots_3_io_debug_p1),
    .io_debug_p2(slots_3_io_debug_p2),
    .io_debug_p3(slots_3_io_debug_p3),
    .io_debug_ppred(slots_3_io_debug_ppred),
    .io_debug_state(slots_3_io_debug_state)
  );
  IssueSlot_16 slots_4 ( // @[issue-unit.scala 157:73]
    .clock(slots_4_clock),
    .reset(slots_4_reset),
    .io_valid(slots_4_io_valid),
    .io_will_be_valid(slots_4_io_will_be_valid),
    .io_request(slots_4_io_request),
    .io_request_hp(slots_4_io_request_hp),
    .io_grant(slots_4_io_grant),
    .io_brupdate_b1_resolve_mask(slots_4_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_4_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_4_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_4_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_4_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_4_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_4_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_4_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_4_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_4_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_4_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_4_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_4_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_4_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_4_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_4_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_4_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_4_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_4_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_4_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_4_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_4_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_4_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_4_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_4_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_4_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_4_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_4_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_4_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_4_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_4_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_4_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_4_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_4_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_4_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_4_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_4_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_4_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_4_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_4_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_4_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_4_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_4_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_4_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_4_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_4_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_4_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_4_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_4_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_4_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_4_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_4_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_4_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_4_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_4_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_4_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_4_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_4_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_4_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_4_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_4_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_4_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_4_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_4_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_4_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_4_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_4_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_4_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_4_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_4_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_4_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_4_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_4_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_4_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_4_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_4_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_4_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_4_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_4_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_4_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_4_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_4_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_4_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_4_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_4_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_4_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_4_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_4_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_4_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_4_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_4_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_4_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_4_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_4_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_4_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_4_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_4_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_4_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_4_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_4_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_4_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_4_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_4_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_4_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_4_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_4_io_brupdate_b2_target_offset),
    .io_kill(slots_4_io_kill),
    .io_clear(slots_4_io_clear),
    .io_ldspec_miss(slots_4_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_4_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_4_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_4_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_4_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_4_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_4_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_4_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_4_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_4_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_4_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_4_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_4_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_4_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_4_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_4_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_4_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_4_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_4_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_4_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_4_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_4_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_4_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_4_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_4_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_4_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_4_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_4_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_4_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_4_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_4_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_4_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_4_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_4_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_4_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_4_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_4_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_4_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_4_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_4_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_4_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_4_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_4_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_4_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_4_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_4_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_4_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_4_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_4_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_4_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_4_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_4_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_4_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_4_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_4_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_4_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_4_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_4_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_4_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_4_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_4_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_4_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_4_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_4_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_4_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_4_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_4_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_4_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_4_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_4_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_4_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_4_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_4_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_4_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_4_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_4_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_4_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_4_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_4_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_4_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_4_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_4_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_4_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_4_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_4_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_4_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_4_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_4_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_4_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_4_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_4_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_4_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_4_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_4_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_4_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_4_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_4_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_4_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_4_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_4_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_4_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_4_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_4_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_4_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_4_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_4_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_4_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_4_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_4_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_4_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_4_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_4_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_4_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_4_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_4_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_4_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_4_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_4_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_4_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_4_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_4_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_4_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_4_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_4_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_4_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_4_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_4_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_4_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_4_io_out_uop_switch),
    .io_out_uop_switch_off(slots_4_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_4_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_4_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_4_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_4_io_out_uop_rflag),
    .io_out_uop_wflag(slots_4_io_out_uop_wflag),
    .io_out_uop_prflag(slots_4_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_4_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_4_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_4_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_4_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_4_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_4_io_out_uop_split_num),
    .io_out_uop_self_index(slots_4_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_4_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_4_io_out_uop_address_num),
    .io_out_uop_uopc(slots_4_io_out_uop_uopc),
    .io_out_uop_inst(slots_4_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_4_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_4_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_4_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_4_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_4_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_4_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_4_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_4_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_4_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_4_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_4_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_4_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_4_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_4_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_4_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_4_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_4_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_4_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_4_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_4_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_4_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_4_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_4_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_4_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_4_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_4_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_4_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_4_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_4_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_4_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_4_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_4_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_4_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_4_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_4_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_4_io_out_uop_pdst),
    .io_out_uop_prs1(slots_4_io_out_uop_prs1),
    .io_out_uop_prs2(slots_4_io_out_uop_prs2),
    .io_out_uop_prs3(slots_4_io_out_uop_prs3),
    .io_out_uop_ppred(slots_4_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_4_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_4_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_4_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_4_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_4_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_4_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_4_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_4_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_4_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_4_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_4_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_4_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_4_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_4_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_4_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_4_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_4_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_4_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_4_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_4_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_4_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_4_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_4_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_4_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_4_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_4_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_4_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_4_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_4_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_4_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_4_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_4_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_4_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_4_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_4_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_4_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_4_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_4_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_4_io_uop_switch),
    .io_uop_switch_off(slots_4_io_uop_switch_off),
    .io_uop_is_unicore(slots_4_io_uop_is_unicore),
    .io_uop_shift(slots_4_io_uop_shift),
    .io_uop_lrs3_rtype(slots_4_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_4_io_uop_rflag),
    .io_uop_wflag(slots_4_io_uop_wflag),
    .io_uop_prflag(slots_4_io_uop_prflag),
    .io_uop_pwflag(slots_4_io_uop_pwflag),
    .io_uop_pflag_busy(slots_4_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_4_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_4_io_uop_op1_sel),
    .io_uop_op2_sel(slots_4_io_uop_op2_sel),
    .io_uop_split_num(slots_4_io_uop_split_num),
    .io_uop_self_index(slots_4_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_4_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_4_io_uop_address_num),
    .io_uop_uopc(slots_4_io_uop_uopc),
    .io_uop_inst(slots_4_io_uop_inst),
    .io_uop_debug_inst(slots_4_io_uop_debug_inst),
    .io_uop_is_rvc(slots_4_io_uop_is_rvc),
    .io_uop_debug_pc(slots_4_io_uop_debug_pc),
    .io_uop_iq_type(slots_4_io_uop_iq_type),
    .io_uop_fu_code(slots_4_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_4_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_4_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_4_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_4_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_4_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_4_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_4_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_4_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_4_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_4_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_4_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_4_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_4_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_4_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_4_io_uop_is_br),
    .io_uop_is_jalr(slots_4_io_uop_is_jalr),
    .io_uop_is_jal(slots_4_io_uop_is_jal),
    .io_uop_is_sfb(slots_4_io_uop_is_sfb),
    .io_uop_br_mask(slots_4_io_uop_br_mask),
    .io_uop_br_tag(slots_4_io_uop_br_tag),
    .io_uop_ftq_idx(slots_4_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_4_io_uop_edge_inst),
    .io_uop_pc_lob(slots_4_io_uop_pc_lob),
    .io_uop_taken(slots_4_io_uop_taken),
    .io_uop_imm_packed(slots_4_io_uop_imm_packed),
    .io_uop_csr_addr(slots_4_io_uop_csr_addr),
    .io_uop_rob_idx(slots_4_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_4_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_4_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_4_io_uop_rxq_idx),
    .io_uop_pdst(slots_4_io_uop_pdst),
    .io_uop_prs1(slots_4_io_uop_prs1),
    .io_uop_prs2(slots_4_io_uop_prs2),
    .io_uop_prs3(slots_4_io_uop_prs3),
    .io_uop_ppred(slots_4_io_uop_ppred),
    .io_uop_prs1_busy(slots_4_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_4_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_4_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_4_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_4_io_uop_stale_pdst),
    .io_uop_exception(slots_4_io_uop_exception),
    .io_uop_exc_cause(slots_4_io_uop_exc_cause),
    .io_uop_bypassable(slots_4_io_uop_bypassable),
    .io_uop_mem_cmd(slots_4_io_uop_mem_cmd),
    .io_uop_mem_size(slots_4_io_uop_mem_size),
    .io_uop_mem_signed(slots_4_io_uop_mem_signed),
    .io_uop_is_fence(slots_4_io_uop_is_fence),
    .io_uop_is_fencei(slots_4_io_uop_is_fencei),
    .io_uop_is_amo(slots_4_io_uop_is_amo),
    .io_uop_uses_ldq(slots_4_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_4_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_4_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_4_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_4_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_4_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_4_io_uop_ldst),
    .io_uop_lrs1(slots_4_io_uop_lrs1),
    .io_uop_lrs2(slots_4_io_uop_lrs2),
    .io_uop_lrs3(slots_4_io_uop_lrs3),
    .io_uop_ldst_val(slots_4_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_4_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_4_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_4_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_4_io_uop_frs3_en),
    .io_uop_fp_val(slots_4_io_uop_fp_val),
    .io_uop_fp_single(slots_4_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_4_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_4_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_4_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_4_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_4_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_4_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_4_io_uop_debug_tsrc),
    .io_debug_p1(slots_4_io_debug_p1),
    .io_debug_p2(slots_4_io_debug_p2),
    .io_debug_p3(slots_4_io_debug_p3),
    .io_debug_ppred(slots_4_io_debug_ppred),
    .io_debug_state(slots_4_io_debug_state)
  );
  IssueSlot_16 slots_5 ( // @[issue-unit.scala 157:73]
    .clock(slots_5_clock),
    .reset(slots_5_reset),
    .io_valid(slots_5_io_valid),
    .io_will_be_valid(slots_5_io_will_be_valid),
    .io_request(slots_5_io_request),
    .io_request_hp(slots_5_io_request_hp),
    .io_grant(slots_5_io_grant),
    .io_brupdate_b1_resolve_mask(slots_5_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_5_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_5_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_5_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_5_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_5_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_5_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_5_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_5_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_5_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_5_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_5_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_5_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_5_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_5_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_5_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_5_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_5_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_5_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_5_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_5_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_5_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_5_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_5_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_5_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_5_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_5_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_5_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_5_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_5_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_5_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_5_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_5_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_5_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_5_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_5_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_5_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_5_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_5_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_5_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_5_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_5_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_5_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_5_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_5_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_5_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_5_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_5_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_5_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_5_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_5_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_5_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_5_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_5_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_5_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_5_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_5_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_5_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_5_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_5_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_5_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_5_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_5_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_5_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_5_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_5_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_5_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_5_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_5_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_5_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_5_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_5_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_5_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_5_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_5_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_5_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_5_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_5_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_5_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_5_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_5_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_5_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_5_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_5_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_5_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_5_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_5_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_5_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_5_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_5_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_5_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_5_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_5_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_5_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_5_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_5_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_5_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_5_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_5_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_5_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_5_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_5_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_5_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_5_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_5_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_5_io_brupdate_b2_target_offset),
    .io_kill(slots_5_io_kill),
    .io_clear(slots_5_io_clear),
    .io_ldspec_miss(slots_5_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_5_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_5_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_5_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_5_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_5_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_5_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_5_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_5_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_5_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_5_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_5_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_5_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_5_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_5_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_5_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_5_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_5_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_5_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_5_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_5_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_5_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_5_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_5_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_5_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_5_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_5_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_5_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_5_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_5_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_5_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_5_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_5_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_5_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_5_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_5_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_5_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_5_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_5_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_5_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_5_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_5_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_5_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_5_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_5_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_5_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_5_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_5_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_5_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_5_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_5_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_5_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_5_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_5_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_5_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_5_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_5_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_5_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_5_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_5_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_5_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_5_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_5_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_5_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_5_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_5_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_5_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_5_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_5_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_5_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_5_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_5_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_5_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_5_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_5_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_5_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_5_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_5_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_5_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_5_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_5_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_5_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_5_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_5_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_5_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_5_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_5_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_5_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_5_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_5_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_5_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_5_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_5_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_5_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_5_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_5_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_5_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_5_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_5_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_5_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_5_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_5_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_5_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_5_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_5_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_5_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_5_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_5_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_5_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_5_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_5_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_5_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_5_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_5_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_5_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_5_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_5_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_5_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_5_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_5_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_5_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_5_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_5_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_5_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_5_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_5_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_5_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_5_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_5_io_out_uop_switch),
    .io_out_uop_switch_off(slots_5_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_5_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_5_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_5_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_5_io_out_uop_rflag),
    .io_out_uop_wflag(slots_5_io_out_uop_wflag),
    .io_out_uop_prflag(slots_5_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_5_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_5_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_5_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_5_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_5_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_5_io_out_uop_split_num),
    .io_out_uop_self_index(slots_5_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_5_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_5_io_out_uop_address_num),
    .io_out_uop_uopc(slots_5_io_out_uop_uopc),
    .io_out_uop_inst(slots_5_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_5_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_5_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_5_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_5_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_5_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_5_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_5_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_5_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_5_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_5_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_5_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_5_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_5_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_5_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_5_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_5_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_5_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_5_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_5_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_5_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_5_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_5_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_5_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_5_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_5_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_5_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_5_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_5_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_5_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_5_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_5_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_5_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_5_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_5_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_5_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_5_io_out_uop_pdst),
    .io_out_uop_prs1(slots_5_io_out_uop_prs1),
    .io_out_uop_prs2(slots_5_io_out_uop_prs2),
    .io_out_uop_prs3(slots_5_io_out_uop_prs3),
    .io_out_uop_ppred(slots_5_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_5_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_5_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_5_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_5_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_5_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_5_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_5_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_5_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_5_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_5_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_5_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_5_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_5_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_5_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_5_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_5_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_5_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_5_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_5_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_5_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_5_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_5_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_5_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_5_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_5_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_5_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_5_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_5_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_5_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_5_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_5_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_5_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_5_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_5_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_5_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_5_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_5_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_5_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_5_io_uop_switch),
    .io_uop_switch_off(slots_5_io_uop_switch_off),
    .io_uop_is_unicore(slots_5_io_uop_is_unicore),
    .io_uop_shift(slots_5_io_uop_shift),
    .io_uop_lrs3_rtype(slots_5_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_5_io_uop_rflag),
    .io_uop_wflag(slots_5_io_uop_wflag),
    .io_uop_prflag(slots_5_io_uop_prflag),
    .io_uop_pwflag(slots_5_io_uop_pwflag),
    .io_uop_pflag_busy(slots_5_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_5_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_5_io_uop_op1_sel),
    .io_uop_op2_sel(slots_5_io_uop_op2_sel),
    .io_uop_split_num(slots_5_io_uop_split_num),
    .io_uop_self_index(slots_5_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_5_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_5_io_uop_address_num),
    .io_uop_uopc(slots_5_io_uop_uopc),
    .io_uop_inst(slots_5_io_uop_inst),
    .io_uop_debug_inst(slots_5_io_uop_debug_inst),
    .io_uop_is_rvc(slots_5_io_uop_is_rvc),
    .io_uop_debug_pc(slots_5_io_uop_debug_pc),
    .io_uop_iq_type(slots_5_io_uop_iq_type),
    .io_uop_fu_code(slots_5_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_5_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_5_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_5_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_5_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_5_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_5_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_5_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_5_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_5_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_5_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_5_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_5_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_5_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_5_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_5_io_uop_is_br),
    .io_uop_is_jalr(slots_5_io_uop_is_jalr),
    .io_uop_is_jal(slots_5_io_uop_is_jal),
    .io_uop_is_sfb(slots_5_io_uop_is_sfb),
    .io_uop_br_mask(slots_5_io_uop_br_mask),
    .io_uop_br_tag(slots_5_io_uop_br_tag),
    .io_uop_ftq_idx(slots_5_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_5_io_uop_edge_inst),
    .io_uop_pc_lob(slots_5_io_uop_pc_lob),
    .io_uop_taken(slots_5_io_uop_taken),
    .io_uop_imm_packed(slots_5_io_uop_imm_packed),
    .io_uop_csr_addr(slots_5_io_uop_csr_addr),
    .io_uop_rob_idx(slots_5_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_5_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_5_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_5_io_uop_rxq_idx),
    .io_uop_pdst(slots_5_io_uop_pdst),
    .io_uop_prs1(slots_5_io_uop_prs1),
    .io_uop_prs2(slots_5_io_uop_prs2),
    .io_uop_prs3(slots_5_io_uop_prs3),
    .io_uop_ppred(slots_5_io_uop_ppred),
    .io_uop_prs1_busy(slots_5_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_5_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_5_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_5_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_5_io_uop_stale_pdst),
    .io_uop_exception(slots_5_io_uop_exception),
    .io_uop_exc_cause(slots_5_io_uop_exc_cause),
    .io_uop_bypassable(slots_5_io_uop_bypassable),
    .io_uop_mem_cmd(slots_5_io_uop_mem_cmd),
    .io_uop_mem_size(slots_5_io_uop_mem_size),
    .io_uop_mem_signed(slots_5_io_uop_mem_signed),
    .io_uop_is_fence(slots_5_io_uop_is_fence),
    .io_uop_is_fencei(slots_5_io_uop_is_fencei),
    .io_uop_is_amo(slots_5_io_uop_is_amo),
    .io_uop_uses_ldq(slots_5_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_5_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_5_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_5_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_5_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_5_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_5_io_uop_ldst),
    .io_uop_lrs1(slots_5_io_uop_lrs1),
    .io_uop_lrs2(slots_5_io_uop_lrs2),
    .io_uop_lrs3(slots_5_io_uop_lrs3),
    .io_uop_ldst_val(slots_5_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_5_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_5_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_5_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_5_io_uop_frs3_en),
    .io_uop_fp_val(slots_5_io_uop_fp_val),
    .io_uop_fp_single(slots_5_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_5_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_5_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_5_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_5_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_5_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_5_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_5_io_uop_debug_tsrc),
    .io_debug_p1(slots_5_io_debug_p1),
    .io_debug_p2(slots_5_io_debug_p2),
    .io_debug_p3(slots_5_io_debug_p3),
    .io_debug_ppred(slots_5_io_debug_ppred),
    .io_debug_state(slots_5_io_debug_state)
  );
  IssueSlot_16 slots_6 ( // @[issue-unit.scala 157:73]
    .clock(slots_6_clock),
    .reset(slots_6_reset),
    .io_valid(slots_6_io_valid),
    .io_will_be_valid(slots_6_io_will_be_valid),
    .io_request(slots_6_io_request),
    .io_request_hp(slots_6_io_request_hp),
    .io_grant(slots_6_io_grant),
    .io_brupdate_b1_resolve_mask(slots_6_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_6_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_6_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_6_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_6_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_6_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_6_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_6_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_6_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_6_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_6_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_6_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_6_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_6_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_6_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_6_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_6_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_6_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_6_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_6_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_6_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_6_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_6_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_6_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_6_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_6_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_6_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_6_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_6_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_6_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_6_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_6_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_6_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_6_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_6_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_6_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_6_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_6_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_6_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_6_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_6_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_6_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_6_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_6_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_6_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_6_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_6_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_6_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_6_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_6_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_6_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_6_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_6_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_6_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_6_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_6_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_6_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_6_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_6_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_6_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_6_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_6_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_6_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_6_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_6_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_6_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_6_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_6_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_6_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_6_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_6_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_6_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_6_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_6_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_6_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_6_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_6_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_6_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_6_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_6_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_6_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_6_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_6_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_6_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_6_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_6_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_6_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_6_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_6_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_6_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_6_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_6_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_6_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_6_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_6_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_6_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_6_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_6_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_6_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_6_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_6_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_6_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_6_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_6_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_6_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_6_io_brupdate_b2_target_offset),
    .io_kill(slots_6_io_kill),
    .io_clear(slots_6_io_clear),
    .io_ldspec_miss(slots_6_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_6_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_6_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_6_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_6_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_6_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_6_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_6_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_6_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_6_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_6_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_6_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_6_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_6_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_6_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_6_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_6_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_6_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_6_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_6_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_6_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_6_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_6_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_6_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_6_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_6_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_6_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_6_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_6_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_6_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_6_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_6_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_6_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_6_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_6_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_6_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_6_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_6_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_6_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_6_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_6_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_6_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_6_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_6_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_6_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_6_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_6_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_6_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_6_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_6_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_6_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_6_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_6_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_6_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_6_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_6_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_6_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_6_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_6_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_6_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_6_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_6_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_6_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_6_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_6_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_6_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_6_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_6_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_6_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_6_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_6_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_6_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_6_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_6_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_6_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_6_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_6_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_6_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_6_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_6_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_6_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_6_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_6_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_6_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_6_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_6_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_6_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_6_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_6_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_6_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_6_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_6_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_6_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_6_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_6_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_6_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_6_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_6_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_6_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_6_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_6_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_6_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_6_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_6_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_6_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_6_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_6_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_6_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_6_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_6_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_6_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_6_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_6_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_6_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_6_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_6_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_6_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_6_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_6_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_6_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_6_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_6_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_6_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_6_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_6_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_6_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_6_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_6_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_6_io_out_uop_switch),
    .io_out_uop_switch_off(slots_6_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_6_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_6_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_6_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_6_io_out_uop_rflag),
    .io_out_uop_wflag(slots_6_io_out_uop_wflag),
    .io_out_uop_prflag(slots_6_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_6_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_6_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_6_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_6_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_6_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_6_io_out_uop_split_num),
    .io_out_uop_self_index(slots_6_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_6_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_6_io_out_uop_address_num),
    .io_out_uop_uopc(slots_6_io_out_uop_uopc),
    .io_out_uop_inst(slots_6_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_6_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_6_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_6_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_6_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_6_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_6_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_6_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_6_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_6_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_6_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_6_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_6_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_6_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_6_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_6_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_6_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_6_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_6_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_6_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_6_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_6_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_6_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_6_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_6_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_6_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_6_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_6_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_6_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_6_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_6_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_6_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_6_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_6_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_6_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_6_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_6_io_out_uop_pdst),
    .io_out_uop_prs1(slots_6_io_out_uop_prs1),
    .io_out_uop_prs2(slots_6_io_out_uop_prs2),
    .io_out_uop_prs3(slots_6_io_out_uop_prs3),
    .io_out_uop_ppred(slots_6_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_6_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_6_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_6_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_6_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_6_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_6_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_6_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_6_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_6_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_6_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_6_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_6_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_6_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_6_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_6_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_6_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_6_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_6_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_6_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_6_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_6_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_6_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_6_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_6_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_6_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_6_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_6_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_6_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_6_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_6_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_6_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_6_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_6_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_6_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_6_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_6_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_6_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_6_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_6_io_uop_switch),
    .io_uop_switch_off(slots_6_io_uop_switch_off),
    .io_uop_is_unicore(slots_6_io_uop_is_unicore),
    .io_uop_shift(slots_6_io_uop_shift),
    .io_uop_lrs3_rtype(slots_6_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_6_io_uop_rflag),
    .io_uop_wflag(slots_6_io_uop_wflag),
    .io_uop_prflag(slots_6_io_uop_prflag),
    .io_uop_pwflag(slots_6_io_uop_pwflag),
    .io_uop_pflag_busy(slots_6_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_6_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_6_io_uop_op1_sel),
    .io_uop_op2_sel(slots_6_io_uop_op2_sel),
    .io_uop_split_num(slots_6_io_uop_split_num),
    .io_uop_self_index(slots_6_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_6_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_6_io_uop_address_num),
    .io_uop_uopc(slots_6_io_uop_uopc),
    .io_uop_inst(slots_6_io_uop_inst),
    .io_uop_debug_inst(slots_6_io_uop_debug_inst),
    .io_uop_is_rvc(slots_6_io_uop_is_rvc),
    .io_uop_debug_pc(slots_6_io_uop_debug_pc),
    .io_uop_iq_type(slots_6_io_uop_iq_type),
    .io_uop_fu_code(slots_6_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_6_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_6_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_6_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_6_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_6_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_6_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_6_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_6_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_6_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_6_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_6_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_6_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_6_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_6_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_6_io_uop_is_br),
    .io_uop_is_jalr(slots_6_io_uop_is_jalr),
    .io_uop_is_jal(slots_6_io_uop_is_jal),
    .io_uop_is_sfb(slots_6_io_uop_is_sfb),
    .io_uop_br_mask(slots_6_io_uop_br_mask),
    .io_uop_br_tag(slots_6_io_uop_br_tag),
    .io_uop_ftq_idx(slots_6_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_6_io_uop_edge_inst),
    .io_uop_pc_lob(slots_6_io_uop_pc_lob),
    .io_uop_taken(slots_6_io_uop_taken),
    .io_uop_imm_packed(slots_6_io_uop_imm_packed),
    .io_uop_csr_addr(slots_6_io_uop_csr_addr),
    .io_uop_rob_idx(slots_6_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_6_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_6_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_6_io_uop_rxq_idx),
    .io_uop_pdst(slots_6_io_uop_pdst),
    .io_uop_prs1(slots_6_io_uop_prs1),
    .io_uop_prs2(slots_6_io_uop_prs2),
    .io_uop_prs3(slots_6_io_uop_prs3),
    .io_uop_ppred(slots_6_io_uop_ppred),
    .io_uop_prs1_busy(slots_6_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_6_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_6_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_6_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_6_io_uop_stale_pdst),
    .io_uop_exception(slots_6_io_uop_exception),
    .io_uop_exc_cause(slots_6_io_uop_exc_cause),
    .io_uop_bypassable(slots_6_io_uop_bypassable),
    .io_uop_mem_cmd(slots_6_io_uop_mem_cmd),
    .io_uop_mem_size(slots_6_io_uop_mem_size),
    .io_uop_mem_signed(slots_6_io_uop_mem_signed),
    .io_uop_is_fence(slots_6_io_uop_is_fence),
    .io_uop_is_fencei(slots_6_io_uop_is_fencei),
    .io_uop_is_amo(slots_6_io_uop_is_amo),
    .io_uop_uses_ldq(slots_6_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_6_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_6_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_6_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_6_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_6_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_6_io_uop_ldst),
    .io_uop_lrs1(slots_6_io_uop_lrs1),
    .io_uop_lrs2(slots_6_io_uop_lrs2),
    .io_uop_lrs3(slots_6_io_uop_lrs3),
    .io_uop_ldst_val(slots_6_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_6_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_6_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_6_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_6_io_uop_frs3_en),
    .io_uop_fp_val(slots_6_io_uop_fp_val),
    .io_uop_fp_single(slots_6_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_6_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_6_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_6_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_6_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_6_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_6_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_6_io_uop_debug_tsrc),
    .io_debug_p1(slots_6_io_debug_p1),
    .io_debug_p2(slots_6_io_debug_p2),
    .io_debug_p3(slots_6_io_debug_p3),
    .io_debug_ppred(slots_6_io_debug_ppred),
    .io_debug_state(slots_6_io_debug_state)
  );
  IssueSlot_16 slots_7 ( // @[issue-unit.scala 157:73]
    .clock(slots_7_clock),
    .reset(slots_7_reset),
    .io_valid(slots_7_io_valid),
    .io_will_be_valid(slots_7_io_will_be_valid),
    .io_request(slots_7_io_request),
    .io_request_hp(slots_7_io_request_hp),
    .io_grant(slots_7_io_grant),
    .io_brupdate_b1_resolve_mask(slots_7_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_7_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_7_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_7_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_7_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_7_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_7_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_7_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_7_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_7_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_7_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_7_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_7_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_7_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_7_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_7_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_7_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_7_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_7_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_7_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_7_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_7_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_7_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_7_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_7_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_7_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_7_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_7_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_7_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_7_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_7_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_7_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_7_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_7_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_7_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_7_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_7_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_7_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_7_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_7_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_7_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_7_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_7_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_7_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_7_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_7_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_7_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_7_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_7_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_7_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_7_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_7_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_7_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_7_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_7_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_7_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_7_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_7_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_7_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_7_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_7_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_7_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_7_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_7_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_7_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_7_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_7_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_7_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_7_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_7_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_7_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_7_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_7_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_7_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_7_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_7_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_7_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_7_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_7_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_7_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_7_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_7_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_7_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_7_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_7_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_7_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_7_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_7_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_7_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_7_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_7_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_7_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_7_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_7_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_7_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_7_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_7_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_7_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_7_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_7_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_7_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_7_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_7_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_7_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_7_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_7_io_brupdate_b2_target_offset),
    .io_kill(slots_7_io_kill),
    .io_clear(slots_7_io_clear),
    .io_ldspec_miss(slots_7_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_7_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_7_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_7_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_7_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_7_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_7_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_7_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_7_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_7_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_7_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_7_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_7_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_7_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_7_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_7_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_7_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_7_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_7_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_7_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_7_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_7_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_7_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_7_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_7_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_7_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_7_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_7_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_7_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_7_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_7_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_7_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_7_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_7_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_7_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_7_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_7_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_7_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_7_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_7_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_7_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_7_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_7_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_7_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_7_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_7_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_7_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_7_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_7_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_7_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_7_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_7_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_7_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_7_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_7_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_7_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_7_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_7_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_7_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_7_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_7_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_7_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_7_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_7_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_7_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_7_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_7_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_7_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_7_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_7_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_7_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_7_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_7_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_7_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_7_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_7_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_7_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_7_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_7_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_7_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_7_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_7_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_7_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_7_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_7_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_7_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_7_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_7_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_7_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_7_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_7_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_7_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_7_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_7_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_7_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_7_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_7_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_7_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_7_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_7_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_7_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_7_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_7_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_7_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_7_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_7_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_7_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_7_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_7_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_7_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_7_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_7_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_7_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_7_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_7_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_7_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_7_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_7_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_7_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_7_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_7_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_7_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_7_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_7_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_7_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_7_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_7_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_7_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_7_io_out_uop_switch),
    .io_out_uop_switch_off(slots_7_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_7_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_7_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_7_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_7_io_out_uop_rflag),
    .io_out_uop_wflag(slots_7_io_out_uop_wflag),
    .io_out_uop_prflag(slots_7_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_7_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_7_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_7_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_7_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_7_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_7_io_out_uop_split_num),
    .io_out_uop_self_index(slots_7_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_7_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_7_io_out_uop_address_num),
    .io_out_uop_uopc(slots_7_io_out_uop_uopc),
    .io_out_uop_inst(slots_7_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_7_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_7_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_7_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_7_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_7_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_7_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_7_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_7_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_7_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_7_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_7_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_7_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_7_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_7_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_7_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_7_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_7_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_7_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_7_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_7_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_7_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_7_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_7_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_7_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_7_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_7_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_7_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_7_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_7_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_7_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_7_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_7_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_7_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_7_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_7_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_7_io_out_uop_pdst),
    .io_out_uop_prs1(slots_7_io_out_uop_prs1),
    .io_out_uop_prs2(slots_7_io_out_uop_prs2),
    .io_out_uop_prs3(slots_7_io_out_uop_prs3),
    .io_out_uop_ppred(slots_7_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_7_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_7_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_7_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_7_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_7_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_7_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_7_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_7_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_7_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_7_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_7_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_7_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_7_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_7_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_7_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_7_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_7_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_7_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_7_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_7_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_7_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_7_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_7_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_7_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_7_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_7_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_7_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_7_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_7_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_7_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_7_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_7_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_7_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_7_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_7_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_7_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_7_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_7_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_7_io_uop_switch),
    .io_uop_switch_off(slots_7_io_uop_switch_off),
    .io_uop_is_unicore(slots_7_io_uop_is_unicore),
    .io_uop_shift(slots_7_io_uop_shift),
    .io_uop_lrs3_rtype(slots_7_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_7_io_uop_rflag),
    .io_uop_wflag(slots_7_io_uop_wflag),
    .io_uop_prflag(slots_7_io_uop_prflag),
    .io_uop_pwflag(slots_7_io_uop_pwflag),
    .io_uop_pflag_busy(slots_7_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_7_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_7_io_uop_op1_sel),
    .io_uop_op2_sel(slots_7_io_uop_op2_sel),
    .io_uop_split_num(slots_7_io_uop_split_num),
    .io_uop_self_index(slots_7_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_7_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_7_io_uop_address_num),
    .io_uop_uopc(slots_7_io_uop_uopc),
    .io_uop_inst(slots_7_io_uop_inst),
    .io_uop_debug_inst(slots_7_io_uop_debug_inst),
    .io_uop_is_rvc(slots_7_io_uop_is_rvc),
    .io_uop_debug_pc(slots_7_io_uop_debug_pc),
    .io_uop_iq_type(slots_7_io_uop_iq_type),
    .io_uop_fu_code(slots_7_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_7_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_7_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_7_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_7_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_7_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_7_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_7_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_7_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_7_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_7_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_7_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_7_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_7_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_7_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_7_io_uop_is_br),
    .io_uop_is_jalr(slots_7_io_uop_is_jalr),
    .io_uop_is_jal(slots_7_io_uop_is_jal),
    .io_uop_is_sfb(slots_7_io_uop_is_sfb),
    .io_uop_br_mask(slots_7_io_uop_br_mask),
    .io_uop_br_tag(slots_7_io_uop_br_tag),
    .io_uop_ftq_idx(slots_7_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_7_io_uop_edge_inst),
    .io_uop_pc_lob(slots_7_io_uop_pc_lob),
    .io_uop_taken(slots_7_io_uop_taken),
    .io_uop_imm_packed(slots_7_io_uop_imm_packed),
    .io_uop_csr_addr(slots_7_io_uop_csr_addr),
    .io_uop_rob_idx(slots_7_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_7_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_7_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_7_io_uop_rxq_idx),
    .io_uop_pdst(slots_7_io_uop_pdst),
    .io_uop_prs1(slots_7_io_uop_prs1),
    .io_uop_prs2(slots_7_io_uop_prs2),
    .io_uop_prs3(slots_7_io_uop_prs3),
    .io_uop_ppred(slots_7_io_uop_ppred),
    .io_uop_prs1_busy(slots_7_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_7_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_7_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_7_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_7_io_uop_stale_pdst),
    .io_uop_exception(slots_7_io_uop_exception),
    .io_uop_exc_cause(slots_7_io_uop_exc_cause),
    .io_uop_bypassable(slots_7_io_uop_bypassable),
    .io_uop_mem_cmd(slots_7_io_uop_mem_cmd),
    .io_uop_mem_size(slots_7_io_uop_mem_size),
    .io_uop_mem_signed(slots_7_io_uop_mem_signed),
    .io_uop_is_fence(slots_7_io_uop_is_fence),
    .io_uop_is_fencei(slots_7_io_uop_is_fencei),
    .io_uop_is_amo(slots_7_io_uop_is_amo),
    .io_uop_uses_ldq(slots_7_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_7_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_7_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_7_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_7_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_7_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_7_io_uop_ldst),
    .io_uop_lrs1(slots_7_io_uop_lrs1),
    .io_uop_lrs2(slots_7_io_uop_lrs2),
    .io_uop_lrs3(slots_7_io_uop_lrs3),
    .io_uop_ldst_val(slots_7_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_7_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_7_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_7_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_7_io_uop_frs3_en),
    .io_uop_fp_val(slots_7_io_uop_fp_val),
    .io_uop_fp_single(slots_7_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_7_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_7_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_7_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_7_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_7_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_7_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_7_io_uop_debug_tsrc),
    .io_debug_p1(slots_7_io_debug_p1),
    .io_debug_p2(slots_7_io_debug_p2),
    .io_debug_p3(slots_7_io_debug_p3),
    .io_debug_ppred(slots_7_io_debug_ppred),
    .io_debug_state(slots_7_io_debug_state)
  );
  IssueSlot_16 slots_8 ( // @[issue-unit.scala 157:73]
    .clock(slots_8_clock),
    .reset(slots_8_reset),
    .io_valid(slots_8_io_valid),
    .io_will_be_valid(slots_8_io_will_be_valid),
    .io_request(slots_8_io_request),
    .io_request_hp(slots_8_io_request_hp),
    .io_grant(slots_8_io_grant),
    .io_brupdate_b1_resolve_mask(slots_8_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_8_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_8_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_8_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_8_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_8_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_8_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_8_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_8_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_8_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_8_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_8_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_8_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_8_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_8_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_8_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_8_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_8_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_8_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_8_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_8_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_8_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_8_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_8_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_8_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_8_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_8_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_8_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_8_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_8_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_8_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_8_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_8_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_8_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_8_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_8_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_8_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_8_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_8_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_8_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_8_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_8_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_8_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_8_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_8_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_8_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_8_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_8_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_8_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_8_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_8_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_8_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_8_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_8_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_8_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_8_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_8_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_8_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_8_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_8_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_8_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_8_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_8_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_8_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_8_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_8_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_8_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_8_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_8_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_8_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_8_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_8_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_8_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_8_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_8_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_8_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_8_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_8_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_8_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_8_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_8_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_8_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_8_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_8_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_8_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_8_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_8_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_8_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_8_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_8_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_8_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_8_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_8_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_8_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_8_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_8_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_8_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_8_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_8_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_8_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_8_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_8_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_8_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_8_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_8_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_8_io_brupdate_b2_target_offset),
    .io_kill(slots_8_io_kill),
    .io_clear(slots_8_io_clear),
    .io_ldspec_miss(slots_8_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_8_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_8_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_8_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_8_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_8_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_8_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_8_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_8_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_8_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_8_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_8_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_8_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_8_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_8_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_8_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_8_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_8_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_8_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_8_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_8_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_8_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_8_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_8_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_8_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_8_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_8_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_8_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_8_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_8_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_8_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_8_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_8_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_8_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_8_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_8_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_8_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_8_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_8_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_8_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_8_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_8_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_8_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_8_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_8_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_8_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_8_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_8_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_8_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_8_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_8_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_8_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_8_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_8_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_8_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_8_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_8_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_8_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_8_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_8_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_8_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_8_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_8_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_8_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_8_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_8_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_8_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_8_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_8_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_8_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_8_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_8_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_8_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_8_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_8_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_8_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_8_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_8_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_8_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_8_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_8_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_8_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_8_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_8_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_8_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_8_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_8_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_8_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_8_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_8_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_8_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_8_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_8_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_8_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_8_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_8_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_8_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_8_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_8_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_8_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_8_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_8_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_8_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_8_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_8_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_8_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_8_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_8_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_8_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_8_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_8_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_8_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_8_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_8_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_8_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_8_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_8_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_8_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_8_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_8_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_8_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_8_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_8_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_8_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_8_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_8_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_8_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_8_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_8_io_out_uop_switch),
    .io_out_uop_switch_off(slots_8_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_8_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_8_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_8_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_8_io_out_uop_rflag),
    .io_out_uop_wflag(slots_8_io_out_uop_wflag),
    .io_out_uop_prflag(slots_8_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_8_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_8_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_8_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_8_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_8_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_8_io_out_uop_split_num),
    .io_out_uop_self_index(slots_8_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_8_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_8_io_out_uop_address_num),
    .io_out_uop_uopc(slots_8_io_out_uop_uopc),
    .io_out_uop_inst(slots_8_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_8_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_8_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_8_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_8_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_8_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_8_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_8_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_8_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_8_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_8_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_8_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_8_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_8_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_8_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_8_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_8_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_8_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_8_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_8_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_8_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_8_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_8_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_8_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_8_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_8_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_8_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_8_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_8_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_8_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_8_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_8_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_8_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_8_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_8_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_8_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_8_io_out_uop_pdst),
    .io_out_uop_prs1(slots_8_io_out_uop_prs1),
    .io_out_uop_prs2(slots_8_io_out_uop_prs2),
    .io_out_uop_prs3(slots_8_io_out_uop_prs3),
    .io_out_uop_ppred(slots_8_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_8_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_8_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_8_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_8_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_8_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_8_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_8_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_8_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_8_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_8_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_8_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_8_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_8_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_8_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_8_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_8_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_8_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_8_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_8_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_8_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_8_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_8_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_8_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_8_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_8_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_8_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_8_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_8_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_8_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_8_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_8_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_8_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_8_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_8_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_8_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_8_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_8_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_8_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_8_io_uop_switch),
    .io_uop_switch_off(slots_8_io_uop_switch_off),
    .io_uop_is_unicore(slots_8_io_uop_is_unicore),
    .io_uop_shift(slots_8_io_uop_shift),
    .io_uop_lrs3_rtype(slots_8_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_8_io_uop_rflag),
    .io_uop_wflag(slots_8_io_uop_wflag),
    .io_uop_prflag(slots_8_io_uop_prflag),
    .io_uop_pwflag(slots_8_io_uop_pwflag),
    .io_uop_pflag_busy(slots_8_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_8_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_8_io_uop_op1_sel),
    .io_uop_op2_sel(slots_8_io_uop_op2_sel),
    .io_uop_split_num(slots_8_io_uop_split_num),
    .io_uop_self_index(slots_8_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_8_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_8_io_uop_address_num),
    .io_uop_uopc(slots_8_io_uop_uopc),
    .io_uop_inst(slots_8_io_uop_inst),
    .io_uop_debug_inst(slots_8_io_uop_debug_inst),
    .io_uop_is_rvc(slots_8_io_uop_is_rvc),
    .io_uop_debug_pc(slots_8_io_uop_debug_pc),
    .io_uop_iq_type(slots_8_io_uop_iq_type),
    .io_uop_fu_code(slots_8_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_8_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_8_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_8_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_8_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_8_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_8_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_8_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_8_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_8_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_8_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_8_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_8_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_8_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_8_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_8_io_uop_is_br),
    .io_uop_is_jalr(slots_8_io_uop_is_jalr),
    .io_uop_is_jal(slots_8_io_uop_is_jal),
    .io_uop_is_sfb(slots_8_io_uop_is_sfb),
    .io_uop_br_mask(slots_8_io_uop_br_mask),
    .io_uop_br_tag(slots_8_io_uop_br_tag),
    .io_uop_ftq_idx(slots_8_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_8_io_uop_edge_inst),
    .io_uop_pc_lob(slots_8_io_uop_pc_lob),
    .io_uop_taken(slots_8_io_uop_taken),
    .io_uop_imm_packed(slots_8_io_uop_imm_packed),
    .io_uop_csr_addr(slots_8_io_uop_csr_addr),
    .io_uop_rob_idx(slots_8_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_8_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_8_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_8_io_uop_rxq_idx),
    .io_uop_pdst(slots_8_io_uop_pdst),
    .io_uop_prs1(slots_8_io_uop_prs1),
    .io_uop_prs2(slots_8_io_uop_prs2),
    .io_uop_prs3(slots_8_io_uop_prs3),
    .io_uop_ppred(slots_8_io_uop_ppred),
    .io_uop_prs1_busy(slots_8_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_8_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_8_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_8_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_8_io_uop_stale_pdst),
    .io_uop_exception(slots_8_io_uop_exception),
    .io_uop_exc_cause(slots_8_io_uop_exc_cause),
    .io_uop_bypassable(slots_8_io_uop_bypassable),
    .io_uop_mem_cmd(slots_8_io_uop_mem_cmd),
    .io_uop_mem_size(slots_8_io_uop_mem_size),
    .io_uop_mem_signed(slots_8_io_uop_mem_signed),
    .io_uop_is_fence(slots_8_io_uop_is_fence),
    .io_uop_is_fencei(slots_8_io_uop_is_fencei),
    .io_uop_is_amo(slots_8_io_uop_is_amo),
    .io_uop_uses_ldq(slots_8_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_8_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_8_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_8_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_8_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_8_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_8_io_uop_ldst),
    .io_uop_lrs1(slots_8_io_uop_lrs1),
    .io_uop_lrs2(slots_8_io_uop_lrs2),
    .io_uop_lrs3(slots_8_io_uop_lrs3),
    .io_uop_ldst_val(slots_8_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_8_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_8_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_8_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_8_io_uop_frs3_en),
    .io_uop_fp_val(slots_8_io_uop_fp_val),
    .io_uop_fp_single(slots_8_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_8_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_8_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_8_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_8_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_8_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_8_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_8_io_uop_debug_tsrc),
    .io_debug_p1(slots_8_io_debug_p1),
    .io_debug_p2(slots_8_io_debug_p2),
    .io_debug_p3(slots_8_io_debug_p3),
    .io_debug_ppred(slots_8_io_debug_ppred),
    .io_debug_state(slots_8_io_debug_state)
  );
  IssueSlot_16 slots_9 ( // @[issue-unit.scala 157:73]
    .clock(slots_9_clock),
    .reset(slots_9_reset),
    .io_valid(slots_9_io_valid),
    .io_will_be_valid(slots_9_io_will_be_valid),
    .io_request(slots_9_io_request),
    .io_request_hp(slots_9_io_request_hp),
    .io_grant(slots_9_io_grant),
    .io_brupdate_b1_resolve_mask(slots_9_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_9_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_9_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_9_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_9_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_9_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_9_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_9_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_9_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_9_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_9_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_9_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_9_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_9_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_9_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_9_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_9_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_9_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_9_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_9_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_9_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_9_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_9_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_9_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_9_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_9_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_9_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_9_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_9_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_9_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_9_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_9_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_9_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_9_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_9_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_9_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_9_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_9_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_9_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_9_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_9_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_9_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_9_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_9_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_9_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_9_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_9_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_9_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_9_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_9_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_9_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_9_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_9_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_9_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_9_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_9_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_9_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_9_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_9_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_9_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_9_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_9_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_9_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_9_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_9_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_9_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_9_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_9_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_9_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_9_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_9_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_9_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_9_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_9_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_9_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_9_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_9_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_9_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_9_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_9_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_9_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_9_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_9_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_9_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_9_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_9_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_9_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_9_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_9_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_9_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_9_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_9_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_9_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_9_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_9_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_9_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_9_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_9_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_9_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_9_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_9_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_9_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_9_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_9_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_9_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_9_io_brupdate_b2_target_offset),
    .io_kill(slots_9_io_kill),
    .io_clear(slots_9_io_clear),
    .io_ldspec_miss(slots_9_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_9_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_9_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_9_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_9_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_9_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_9_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_9_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_9_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_9_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_9_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_9_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_9_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_9_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_9_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_9_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_9_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_9_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_9_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_9_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_9_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_9_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_9_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_9_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_9_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_9_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_9_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_9_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_9_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_9_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_9_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_9_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_9_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_9_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_9_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_9_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_9_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_9_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_9_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_9_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_9_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_9_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_9_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_9_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_9_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_9_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_9_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_9_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_9_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_9_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_9_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_9_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_9_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_9_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_9_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_9_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_9_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_9_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_9_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_9_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_9_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_9_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_9_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_9_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_9_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_9_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_9_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_9_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_9_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_9_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_9_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_9_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_9_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_9_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_9_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_9_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_9_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_9_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_9_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_9_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_9_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_9_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_9_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_9_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_9_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_9_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_9_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_9_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_9_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_9_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_9_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_9_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_9_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_9_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_9_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_9_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_9_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_9_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_9_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_9_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_9_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_9_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_9_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_9_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_9_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_9_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_9_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_9_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_9_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_9_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_9_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_9_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_9_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_9_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_9_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_9_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_9_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_9_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_9_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_9_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_9_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_9_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_9_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_9_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_9_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_9_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_9_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_9_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_9_io_out_uop_switch),
    .io_out_uop_switch_off(slots_9_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_9_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_9_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_9_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_9_io_out_uop_rflag),
    .io_out_uop_wflag(slots_9_io_out_uop_wflag),
    .io_out_uop_prflag(slots_9_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_9_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_9_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_9_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_9_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_9_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_9_io_out_uop_split_num),
    .io_out_uop_self_index(slots_9_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_9_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_9_io_out_uop_address_num),
    .io_out_uop_uopc(slots_9_io_out_uop_uopc),
    .io_out_uop_inst(slots_9_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_9_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_9_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_9_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_9_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_9_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_9_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_9_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_9_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_9_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_9_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_9_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_9_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_9_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_9_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_9_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_9_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_9_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_9_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_9_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_9_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_9_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_9_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_9_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_9_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_9_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_9_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_9_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_9_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_9_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_9_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_9_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_9_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_9_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_9_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_9_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_9_io_out_uop_pdst),
    .io_out_uop_prs1(slots_9_io_out_uop_prs1),
    .io_out_uop_prs2(slots_9_io_out_uop_prs2),
    .io_out_uop_prs3(slots_9_io_out_uop_prs3),
    .io_out_uop_ppred(slots_9_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_9_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_9_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_9_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_9_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_9_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_9_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_9_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_9_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_9_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_9_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_9_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_9_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_9_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_9_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_9_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_9_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_9_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_9_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_9_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_9_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_9_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_9_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_9_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_9_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_9_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_9_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_9_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_9_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_9_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_9_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_9_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_9_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_9_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_9_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_9_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_9_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_9_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_9_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_9_io_uop_switch),
    .io_uop_switch_off(slots_9_io_uop_switch_off),
    .io_uop_is_unicore(slots_9_io_uop_is_unicore),
    .io_uop_shift(slots_9_io_uop_shift),
    .io_uop_lrs3_rtype(slots_9_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_9_io_uop_rflag),
    .io_uop_wflag(slots_9_io_uop_wflag),
    .io_uop_prflag(slots_9_io_uop_prflag),
    .io_uop_pwflag(slots_9_io_uop_pwflag),
    .io_uop_pflag_busy(slots_9_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_9_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_9_io_uop_op1_sel),
    .io_uop_op2_sel(slots_9_io_uop_op2_sel),
    .io_uop_split_num(slots_9_io_uop_split_num),
    .io_uop_self_index(slots_9_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_9_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_9_io_uop_address_num),
    .io_uop_uopc(slots_9_io_uop_uopc),
    .io_uop_inst(slots_9_io_uop_inst),
    .io_uop_debug_inst(slots_9_io_uop_debug_inst),
    .io_uop_is_rvc(slots_9_io_uop_is_rvc),
    .io_uop_debug_pc(slots_9_io_uop_debug_pc),
    .io_uop_iq_type(slots_9_io_uop_iq_type),
    .io_uop_fu_code(slots_9_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_9_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_9_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_9_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_9_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_9_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_9_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_9_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_9_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_9_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_9_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_9_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_9_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_9_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_9_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_9_io_uop_is_br),
    .io_uop_is_jalr(slots_9_io_uop_is_jalr),
    .io_uop_is_jal(slots_9_io_uop_is_jal),
    .io_uop_is_sfb(slots_9_io_uop_is_sfb),
    .io_uop_br_mask(slots_9_io_uop_br_mask),
    .io_uop_br_tag(slots_9_io_uop_br_tag),
    .io_uop_ftq_idx(slots_9_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_9_io_uop_edge_inst),
    .io_uop_pc_lob(slots_9_io_uop_pc_lob),
    .io_uop_taken(slots_9_io_uop_taken),
    .io_uop_imm_packed(slots_9_io_uop_imm_packed),
    .io_uop_csr_addr(slots_9_io_uop_csr_addr),
    .io_uop_rob_idx(slots_9_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_9_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_9_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_9_io_uop_rxq_idx),
    .io_uop_pdst(slots_9_io_uop_pdst),
    .io_uop_prs1(slots_9_io_uop_prs1),
    .io_uop_prs2(slots_9_io_uop_prs2),
    .io_uop_prs3(slots_9_io_uop_prs3),
    .io_uop_ppred(slots_9_io_uop_ppred),
    .io_uop_prs1_busy(slots_9_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_9_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_9_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_9_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_9_io_uop_stale_pdst),
    .io_uop_exception(slots_9_io_uop_exception),
    .io_uop_exc_cause(slots_9_io_uop_exc_cause),
    .io_uop_bypassable(slots_9_io_uop_bypassable),
    .io_uop_mem_cmd(slots_9_io_uop_mem_cmd),
    .io_uop_mem_size(slots_9_io_uop_mem_size),
    .io_uop_mem_signed(slots_9_io_uop_mem_signed),
    .io_uop_is_fence(slots_9_io_uop_is_fence),
    .io_uop_is_fencei(slots_9_io_uop_is_fencei),
    .io_uop_is_amo(slots_9_io_uop_is_amo),
    .io_uop_uses_ldq(slots_9_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_9_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_9_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_9_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_9_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_9_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_9_io_uop_ldst),
    .io_uop_lrs1(slots_9_io_uop_lrs1),
    .io_uop_lrs2(slots_9_io_uop_lrs2),
    .io_uop_lrs3(slots_9_io_uop_lrs3),
    .io_uop_ldst_val(slots_9_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_9_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_9_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_9_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_9_io_uop_frs3_en),
    .io_uop_fp_val(slots_9_io_uop_fp_val),
    .io_uop_fp_single(slots_9_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_9_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_9_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_9_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_9_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_9_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_9_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_9_io_uop_debug_tsrc),
    .io_debug_p1(slots_9_io_debug_p1),
    .io_debug_p2(slots_9_io_debug_p2),
    .io_debug_p3(slots_9_io_debug_p3),
    .io_debug_ppred(slots_9_io_debug_ppred),
    .io_debug_state(slots_9_io_debug_state)
  );
  IssueSlot_16 slots_10 ( // @[issue-unit.scala 157:73]
    .clock(slots_10_clock),
    .reset(slots_10_reset),
    .io_valid(slots_10_io_valid),
    .io_will_be_valid(slots_10_io_will_be_valid),
    .io_request(slots_10_io_request),
    .io_request_hp(slots_10_io_request_hp),
    .io_grant(slots_10_io_grant),
    .io_brupdate_b1_resolve_mask(slots_10_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_10_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_10_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_10_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_10_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_10_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_10_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_10_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_10_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_10_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_10_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_10_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_10_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_10_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_10_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_10_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_10_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_10_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_10_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_10_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_10_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_10_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_10_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_10_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_10_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_10_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_10_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_10_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_10_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_10_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_10_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_10_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_10_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_10_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_10_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_10_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_10_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_10_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_10_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_10_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_10_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_10_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_10_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_10_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_10_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_10_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_10_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_10_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_10_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_10_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_10_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_10_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_10_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_10_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_10_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_10_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_10_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_10_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_10_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_10_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_10_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_10_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_10_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_10_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_10_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_10_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_10_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_10_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_10_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_10_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_10_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_10_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_10_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_10_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_10_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_10_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_10_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_10_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_10_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_10_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_10_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_10_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_10_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_10_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_10_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_10_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_10_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_10_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_10_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_10_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_10_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_10_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_10_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_10_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_10_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_10_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_10_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_10_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_10_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_10_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_10_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_10_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_10_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_10_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_10_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_10_io_brupdate_b2_target_offset),
    .io_kill(slots_10_io_kill),
    .io_clear(slots_10_io_clear),
    .io_ldspec_miss(slots_10_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_10_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_10_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_10_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_10_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_10_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_10_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_10_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_10_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_10_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_10_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_10_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_10_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_10_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_10_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_10_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_10_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_10_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_10_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_10_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_10_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_10_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_10_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_10_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_10_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_10_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_10_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_10_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_10_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_10_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_10_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_10_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_10_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_10_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_10_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_10_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_10_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_10_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_10_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_10_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_10_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_10_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_10_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_10_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_10_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_10_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_10_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_10_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_10_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_10_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_10_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_10_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_10_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_10_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_10_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_10_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_10_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_10_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_10_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_10_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_10_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_10_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_10_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_10_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_10_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_10_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_10_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_10_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_10_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_10_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_10_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_10_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_10_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_10_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_10_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_10_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_10_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_10_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_10_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_10_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_10_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_10_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_10_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_10_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_10_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_10_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_10_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_10_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_10_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_10_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_10_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_10_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_10_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_10_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_10_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_10_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_10_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_10_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_10_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_10_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_10_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_10_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_10_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_10_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_10_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_10_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_10_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_10_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_10_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_10_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_10_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_10_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_10_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_10_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_10_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_10_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_10_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_10_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_10_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_10_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_10_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_10_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_10_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_10_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_10_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_10_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_10_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_10_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_10_io_out_uop_switch),
    .io_out_uop_switch_off(slots_10_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_10_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_10_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_10_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_10_io_out_uop_rflag),
    .io_out_uop_wflag(slots_10_io_out_uop_wflag),
    .io_out_uop_prflag(slots_10_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_10_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_10_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_10_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_10_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_10_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_10_io_out_uop_split_num),
    .io_out_uop_self_index(slots_10_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_10_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_10_io_out_uop_address_num),
    .io_out_uop_uopc(slots_10_io_out_uop_uopc),
    .io_out_uop_inst(slots_10_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_10_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_10_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_10_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_10_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_10_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_10_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_10_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_10_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_10_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_10_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_10_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_10_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_10_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_10_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_10_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_10_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_10_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_10_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_10_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_10_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_10_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_10_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_10_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_10_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_10_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_10_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_10_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_10_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_10_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_10_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_10_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_10_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_10_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_10_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_10_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_10_io_out_uop_pdst),
    .io_out_uop_prs1(slots_10_io_out_uop_prs1),
    .io_out_uop_prs2(slots_10_io_out_uop_prs2),
    .io_out_uop_prs3(slots_10_io_out_uop_prs3),
    .io_out_uop_ppred(slots_10_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_10_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_10_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_10_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_10_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_10_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_10_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_10_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_10_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_10_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_10_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_10_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_10_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_10_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_10_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_10_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_10_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_10_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_10_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_10_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_10_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_10_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_10_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_10_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_10_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_10_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_10_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_10_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_10_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_10_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_10_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_10_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_10_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_10_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_10_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_10_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_10_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_10_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_10_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_10_io_uop_switch),
    .io_uop_switch_off(slots_10_io_uop_switch_off),
    .io_uop_is_unicore(slots_10_io_uop_is_unicore),
    .io_uop_shift(slots_10_io_uop_shift),
    .io_uop_lrs3_rtype(slots_10_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_10_io_uop_rflag),
    .io_uop_wflag(slots_10_io_uop_wflag),
    .io_uop_prflag(slots_10_io_uop_prflag),
    .io_uop_pwflag(slots_10_io_uop_pwflag),
    .io_uop_pflag_busy(slots_10_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_10_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_10_io_uop_op1_sel),
    .io_uop_op2_sel(slots_10_io_uop_op2_sel),
    .io_uop_split_num(slots_10_io_uop_split_num),
    .io_uop_self_index(slots_10_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_10_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_10_io_uop_address_num),
    .io_uop_uopc(slots_10_io_uop_uopc),
    .io_uop_inst(slots_10_io_uop_inst),
    .io_uop_debug_inst(slots_10_io_uop_debug_inst),
    .io_uop_is_rvc(slots_10_io_uop_is_rvc),
    .io_uop_debug_pc(slots_10_io_uop_debug_pc),
    .io_uop_iq_type(slots_10_io_uop_iq_type),
    .io_uop_fu_code(slots_10_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_10_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_10_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_10_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_10_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_10_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_10_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_10_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_10_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_10_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_10_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_10_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_10_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_10_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_10_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_10_io_uop_is_br),
    .io_uop_is_jalr(slots_10_io_uop_is_jalr),
    .io_uop_is_jal(slots_10_io_uop_is_jal),
    .io_uop_is_sfb(slots_10_io_uop_is_sfb),
    .io_uop_br_mask(slots_10_io_uop_br_mask),
    .io_uop_br_tag(slots_10_io_uop_br_tag),
    .io_uop_ftq_idx(slots_10_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_10_io_uop_edge_inst),
    .io_uop_pc_lob(slots_10_io_uop_pc_lob),
    .io_uop_taken(slots_10_io_uop_taken),
    .io_uop_imm_packed(slots_10_io_uop_imm_packed),
    .io_uop_csr_addr(slots_10_io_uop_csr_addr),
    .io_uop_rob_idx(slots_10_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_10_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_10_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_10_io_uop_rxq_idx),
    .io_uop_pdst(slots_10_io_uop_pdst),
    .io_uop_prs1(slots_10_io_uop_prs1),
    .io_uop_prs2(slots_10_io_uop_prs2),
    .io_uop_prs3(slots_10_io_uop_prs3),
    .io_uop_ppred(slots_10_io_uop_ppred),
    .io_uop_prs1_busy(slots_10_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_10_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_10_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_10_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_10_io_uop_stale_pdst),
    .io_uop_exception(slots_10_io_uop_exception),
    .io_uop_exc_cause(slots_10_io_uop_exc_cause),
    .io_uop_bypassable(slots_10_io_uop_bypassable),
    .io_uop_mem_cmd(slots_10_io_uop_mem_cmd),
    .io_uop_mem_size(slots_10_io_uop_mem_size),
    .io_uop_mem_signed(slots_10_io_uop_mem_signed),
    .io_uop_is_fence(slots_10_io_uop_is_fence),
    .io_uop_is_fencei(slots_10_io_uop_is_fencei),
    .io_uop_is_amo(slots_10_io_uop_is_amo),
    .io_uop_uses_ldq(slots_10_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_10_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_10_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_10_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_10_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_10_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_10_io_uop_ldst),
    .io_uop_lrs1(slots_10_io_uop_lrs1),
    .io_uop_lrs2(slots_10_io_uop_lrs2),
    .io_uop_lrs3(slots_10_io_uop_lrs3),
    .io_uop_ldst_val(slots_10_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_10_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_10_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_10_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_10_io_uop_frs3_en),
    .io_uop_fp_val(slots_10_io_uop_fp_val),
    .io_uop_fp_single(slots_10_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_10_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_10_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_10_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_10_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_10_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_10_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_10_io_uop_debug_tsrc),
    .io_debug_p1(slots_10_io_debug_p1),
    .io_debug_p2(slots_10_io_debug_p2),
    .io_debug_p3(slots_10_io_debug_p3),
    .io_debug_ppred(slots_10_io_debug_ppred),
    .io_debug_state(slots_10_io_debug_state)
  );
  IssueSlot_16 slots_11 ( // @[issue-unit.scala 157:73]
    .clock(slots_11_clock),
    .reset(slots_11_reset),
    .io_valid(slots_11_io_valid),
    .io_will_be_valid(slots_11_io_will_be_valid),
    .io_request(slots_11_io_request),
    .io_request_hp(slots_11_io_request_hp),
    .io_grant(slots_11_io_grant),
    .io_brupdate_b1_resolve_mask(slots_11_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_11_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_11_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_11_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_11_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_11_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_11_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_11_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_11_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_11_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_11_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_11_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_11_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_11_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_11_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_11_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_11_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_11_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_11_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_11_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_11_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_11_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_11_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_11_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_11_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_11_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_11_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_11_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_11_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_11_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_11_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_11_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_11_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_11_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_11_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_11_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_11_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_11_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_11_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_11_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_11_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_11_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_11_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_11_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_11_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_11_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_11_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_11_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_11_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_11_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_11_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_11_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_11_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_11_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_11_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_11_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_11_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_11_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_11_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_11_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_11_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_11_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_11_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_11_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_11_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_11_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_11_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_11_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_11_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_11_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_11_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_11_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_11_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_11_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_11_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_11_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_11_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_11_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_11_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_11_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_11_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_11_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_11_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_11_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_11_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_11_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_11_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_11_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_11_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_11_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_11_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_11_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_11_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_11_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_11_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_11_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_11_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_11_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_11_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_11_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_11_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_11_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_11_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_11_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_11_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_11_io_brupdate_b2_target_offset),
    .io_kill(slots_11_io_kill),
    .io_clear(slots_11_io_clear),
    .io_ldspec_miss(slots_11_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_11_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_11_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_11_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_11_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_11_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_11_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_11_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_11_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_11_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_11_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_11_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_11_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_11_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_11_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_11_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_11_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_11_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_11_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_11_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_11_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_11_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_11_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_11_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_11_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_11_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_11_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_11_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_11_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_11_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_11_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_11_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_11_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_11_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_11_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_11_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_11_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_11_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_11_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_11_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_11_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_11_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_11_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_11_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_11_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_11_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_11_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_11_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_11_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_11_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_11_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_11_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_11_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_11_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_11_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_11_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_11_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_11_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_11_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_11_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_11_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_11_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_11_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_11_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_11_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_11_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_11_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_11_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_11_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_11_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_11_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_11_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_11_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_11_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_11_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_11_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_11_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_11_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_11_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_11_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_11_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_11_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_11_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_11_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_11_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_11_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_11_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_11_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_11_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_11_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_11_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_11_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_11_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_11_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_11_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_11_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_11_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_11_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_11_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_11_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_11_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_11_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_11_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_11_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_11_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_11_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_11_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_11_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_11_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_11_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_11_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_11_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_11_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_11_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_11_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_11_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_11_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_11_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_11_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_11_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_11_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_11_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_11_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_11_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_11_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_11_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_11_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_11_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_11_io_out_uop_switch),
    .io_out_uop_switch_off(slots_11_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_11_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_11_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_11_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_11_io_out_uop_rflag),
    .io_out_uop_wflag(slots_11_io_out_uop_wflag),
    .io_out_uop_prflag(slots_11_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_11_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_11_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_11_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_11_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_11_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_11_io_out_uop_split_num),
    .io_out_uop_self_index(slots_11_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_11_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_11_io_out_uop_address_num),
    .io_out_uop_uopc(slots_11_io_out_uop_uopc),
    .io_out_uop_inst(slots_11_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_11_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_11_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_11_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_11_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_11_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_11_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_11_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_11_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_11_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_11_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_11_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_11_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_11_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_11_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_11_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_11_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_11_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_11_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_11_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_11_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_11_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_11_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_11_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_11_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_11_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_11_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_11_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_11_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_11_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_11_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_11_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_11_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_11_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_11_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_11_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_11_io_out_uop_pdst),
    .io_out_uop_prs1(slots_11_io_out_uop_prs1),
    .io_out_uop_prs2(slots_11_io_out_uop_prs2),
    .io_out_uop_prs3(slots_11_io_out_uop_prs3),
    .io_out_uop_ppred(slots_11_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_11_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_11_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_11_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_11_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_11_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_11_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_11_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_11_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_11_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_11_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_11_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_11_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_11_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_11_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_11_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_11_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_11_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_11_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_11_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_11_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_11_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_11_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_11_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_11_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_11_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_11_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_11_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_11_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_11_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_11_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_11_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_11_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_11_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_11_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_11_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_11_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_11_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_11_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_11_io_uop_switch),
    .io_uop_switch_off(slots_11_io_uop_switch_off),
    .io_uop_is_unicore(slots_11_io_uop_is_unicore),
    .io_uop_shift(slots_11_io_uop_shift),
    .io_uop_lrs3_rtype(slots_11_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_11_io_uop_rflag),
    .io_uop_wflag(slots_11_io_uop_wflag),
    .io_uop_prflag(slots_11_io_uop_prflag),
    .io_uop_pwflag(slots_11_io_uop_pwflag),
    .io_uop_pflag_busy(slots_11_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_11_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_11_io_uop_op1_sel),
    .io_uop_op2_sel(slots_11_io_uop_op2_sel),
    .io_uop_split_num(slots_11_io_uop_split_num),
    .io_uop_self_index(slots_11_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_11_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_11_io_uop_address_num),
    .io_uop_uopc(slots_11_io_uop_uopc),
    .io_uop_inst(slots_11_io_uop_inst),
    .io_uop_debug_inst(slots_11_io_uop_debug_inst),
    .io_uop_is_rvc(slots_11_io_uop_is_rvc),
    .io_uop_debug_pc(slots_11_io_uop_debug_pc),
    .io_uop_iq_type(slots_11_io_uop_iq_type),
    .io_uop_fu_code(slots_11_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_11_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_11_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_11_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_11_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_11_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_11_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_11_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_11_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_11_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_11_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_11_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_11_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_11_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_11_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_11_io_uop_is_br),
    .io_uop_is_jalr(slots_11_io_uop_is_jalr),
    .io_uop_is_jal(slots_11_io_uop_is_jal),
    .io_uop_is_sfb(slots_11_io_uop_is_sfb),
    .io_uop_br_mask(slots_11_io_uop_br_mask),
    .io_uop_br_tag(slots_11_io_uop_br_tag),
    .io_uop_ftq_idx(slots_11_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_11_io_uop_edge_inst),
    .io_uop_pc_lob(slots_11_io_uop_pc_lob),
    .io_uop_taken(slots_11_io_uop_taken),
    .io_uop_imm_packed(slots_11_io_uop_imm_packed),
    .io_uop_csr_addr(slots_11_io_uop_csr_addr),
    .io_uop_rob_idx(slots_11_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_11_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_11_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_11_io_uop_rxq_idx),
    .io_uop_pdst(slots_11_io_uop_pdst),
    .io_uop_prs1(slots_11_io_uop_prs1),
    .io_uop_prs2(slots_11_io_uop_prs2),
    .io_uop_prs3(slots_11_io_uop_prs3),
    .io_uop_ppred(slots_11_io_uop_ppred),
    .io_uop_prs1_busy(slots_11_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_11_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_11_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_11_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_11_io_uop_stale_pdst),
    .io_uop_exception(slots_11_io_uop_exception),
    .io_uop_exc_cause(slots_11_io_uop_exc_cause),
    .io_uop_bypassable(slots_11_io_uop_bypassable),
    .io_uop_mem_cmd(slots_11_io_uop_mem_cmd),
    .io_uop_mem_size(slots_11_io_uop_mem_size),
    .io_uop_mem_signed(slots_11_io_uop_mem_signed),
    .io_uop_is_fence(slots_11_io_uop_is_fence),
    .io_uop_is_fencei(slots_11_io_uop_is_fencei),
    .io_uop_is_amo(slots_11_io_uop_is_amo),
    .io_uop_uses_ldq(slots_11_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_11_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_11_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_11_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_11_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_11_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_11_io_uop_ldst),
    .io_uop_lrs1(slots_11_io_uop_lrs1),
    .io_uop_lrs2(slots_11_io_uop_lrs2),
    .io_uop_lrs3(slots_11_io_uop_lrs3),
    .io_uop_ldst_val(slots_11_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_11_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_11_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_11_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_11_io_uop_frs3_en),
    .io_uop_fp_val(slots_11_io_uop_fp_val),
    .io_uop_fp_single(slots_11_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_11_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_11_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_11_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_11_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_11_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_11_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_11_io_uop_debug_tsrc),
    .io_debug_p1(slots_11_io_debug_p1),
    .io_debug_p2(slots_11_io_debug_p2),
    .io_debug_p3(slots_11_io_debug_p3),
    .io_debug_ppred(slots_11_io_debug_ppred),
    .io_debug_state(slots_11_io_debug_state)
  );
  IssueSlot_16 slots_12 ( // @[issue-unit.scala 157:73]
    .clock(slots_12_clock),
    .reset(slots_12_reset),
    .io_valid(slots_12_io_valid),
    .io_will_be_valid(slots_12_io_will_be_valid),
    .io_request(slots_12_io_request),
    .io_request_hp(slots_12_io_request_hp),
    .io_grant(slots_12_io_grant),
    .io_brupdate_b1_resolve_mask(slots_12_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_12_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_12_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_12_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_12_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_12_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_12_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_12_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_12_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_12_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_12_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_12_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_12_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_12_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_12_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_12_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_12_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_12_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_12_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_12_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_12_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_12_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_12_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_12_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_12_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_12_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_12_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_12_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_12_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_12_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_12_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_12_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_12_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_12_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_12_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_12_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_12_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_12_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_12_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_12_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_12_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_12_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_12_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_12_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_12_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_12_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_12_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_12_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_12_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_12_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_12_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_12_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_12_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_12_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_12_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_12_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_12_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_12_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_12_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_12_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_12_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_12_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_12_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_12_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_12_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_12_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_12_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_12_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_12_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_12_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_12_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_12_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_12_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_12_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_12_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_12_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_12_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_12_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_12_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_12_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_12_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_12_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_12_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_12_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_12_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_12_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_12_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_12_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_12_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_12_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_12_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_12_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_12_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_12_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_12_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_12_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_12_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_12_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_12_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_12_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_12_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_12_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_12_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_12_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_12_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_12_io_brupdate_b2_target_offset),
    .io_kill(slots_12_io_kill),
    .io_clear(slots_12_io_clear),
    .io_ldspec_miss(slots_12_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_12_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_12_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_12_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_12_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_12_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_12_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_12_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_12_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_12_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_12_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_12_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_12_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_12_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_12_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_12_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_12_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_12_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_12_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_12_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_12_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_12_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_12_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_12_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_12_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_12_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_12_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_12_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_12_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_12_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_12_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_12_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_12_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_12_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_12_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_12_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_12_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_12_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_12_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_12_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_12_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_12_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_12_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_12_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_12_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_12_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_12_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_12_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_12_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_12_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_12_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_12_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_12_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_12_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_12_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_12_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_12_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_12_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_12_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_12_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_12_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_12_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_12_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_12_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_12_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_12_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_12_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_12_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_12_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_12_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_12_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_12_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_12_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_12_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_12_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_12_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_12_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_12_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_12_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_12_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_12_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_12_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_12_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_12_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_12_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_12_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_12_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_12_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_12_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_12_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_12_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_12_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_12_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_12_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_12_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_12_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_12_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_12_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_12_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_12_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_12_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_12_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_12_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_12_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_12_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_12_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_12_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_12_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_12_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_12_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_12_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_12_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_12_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_12_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_12_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_12_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_12_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_12_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_12_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_12_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_12_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_12_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_12_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_12_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_12_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_12_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_12_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_12_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_12_io_out_uop_switch),
    .io_out_uop_switch_off(slots_12_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_12_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_12_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_12_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_12_io_out_uop_rflag),
    .io_out_uop_wflag(slots_12_io_out_uop_wflag),
    .io_out_uop_prflag(slots_12_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_12_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_12_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_12_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_12_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_12_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_12_io_out_uop_split_num),
    .io_out_uop_self_index(slots_12_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_12_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_12_io_out_uop_address_num),
    .io_out_uop_uopc(slots_12_io_out_uop_uopc),
    .io_out_uop_inst(slots_12_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_12_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_12_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_12_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_12_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_12_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_12_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_12_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_12_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_12_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_12_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_12_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_12_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_12_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_12_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_12_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_12_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_12_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_12_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_12_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_12_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_12_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_12_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_12_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_12_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_12_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_12_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_12_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_12_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_12_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_12_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_12_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_12_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_12_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_12_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_12_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_12_io_out_uop_pdst),
    .io_out_uop_prs1(slots_12_io_out_uop_prs1),
    .io_out_uop_prs2(slots_12_io_out_uop_prs2),
    .io_out_uop_prs3(slots_12_io_out_uop_prs3),
    .io_out_uop_ppred(slots_12_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_12_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_12_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_12_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_12_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_12_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_12_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_12_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_12_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_12_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_12_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_12_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_12_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_12_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_12_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_12_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_12_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_12_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_12_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_12_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_12_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_12_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_12_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_12_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_12_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_12_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_12_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_12_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_12_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_12_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_12_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_12_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_12_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_12_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_12_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_12_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_12_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_12_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_12_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_12_io_uop_switch),
    .io_uop_switch_off(slots_12_io_uop_switch_off),
    .io_uop_is_unicore(slots_12_io_uop_is_unicore),
    .io_uop_shift(slots_12_io_uop_shift),
    .io_uop_lrs3_rtype(slots_12_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_12_io_uop_rflag),
    .io_uop_wflag(slots_12_io_uop_wflag),
    .io_uop_prflag(slots_12_io_uop_prflag),
    .io_uop_pwflag(slots_12_io_uop_pwflag),
    .io_uop_pflag_busy(slots_12_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_12_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_12_io_uop_op1_sel),
    .io_uop_op2_sel(slots_12_io_uop_op2_sel),
    .io_uop_split_num(slots_12_io_uop_split_num),
    .io_uop_self_index(slots_12_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_12_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_12_io_uop_address_num),
    .io_uop_uopc(slots_12_io_uop_uopc),
    .io_uop_inst(slots_12_io_uop_inst),
    .io_uop_debug_inst(slots_12_io_uop_debug_inst),
    .io_uop_is_rvc(slots_12_io_uop_is_rvc),
    .io_uop_debug_pc(slots_12_io_uop_debug_pc),
    .io_uop_iq_type(slots_12_io_uop_iq_type),
    .io_uop_fu_code(slots_12_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_12_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_12_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_12_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_12_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_12_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_12_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_12_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_12_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_12_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_12_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_12_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_12_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_12_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_12_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_12_io_uop_is_br),
    .io_uop_is_jalr(slots_12_io_uop_is_jalr),
    .io_uop_is_jal(slots_12_io_uop_is_jal),
    .io_uop_is_sfb(slots_12_io_uop_is_sfb),
    .io_uop_br_mask(slots_12_io_uop_br_mask),
    .io_uop_br_tag(slots_12_io_uop_br_tag),
    .io_uop_ftq_idx(slots_12_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_12_io_uop_edge_inst),
    .io_uop_pc_lob(slots_12_io_uop_pc_lob),
    .io_uop_taken(slots_12_io_uop_taken),
    .io_uop_imm_packed(slots_12_io_uop_imm_packed),
    .io_uop_csr_addr(slots_12_io_uop_csr_addr),
    .io_uop_rob_idx(slots_12_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_12_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_12_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_12_io_uop_rxq_idx),
    .io_uop_pdst(slots_12_io_uop_pdst),
    .io_uop_prs1(slots_12_io_uop_prs1),
    .io_uop_prs2(slots_12_io_uop_prs2),
    .io_uop_prs3(slots_12_io_uop_prs3),
    .io_uop_ppred(slots_12_io_uop_ppred),
    .io_uop_prs1_busy(slots_12_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_12_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_12_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_12_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_12_io_uop_stale_pdst),
    .io_uop_exception(slots_12_io_uop_exception),
    .io_uop_exc_cause(slots_12_io_uop_exc_cause),
    .io_uop_bypassable(slots_12_io_uop_bypassable),
    .io_uop_mem_cmd(slots_12_io_uop_mem_cmd),
    .io_uop_mem_size(slots_12_io_uop_mem_size),
    .io_uop_mem_signed(slots_12_io_uop_mem_signed),
    .io_uop_is_fence(slots_12_io_uop_is_fence),
    .io_uop_is_fencei(slots_12_io_uop_is_fencei),
    .io_uop_is_amo(slots_12_io_uop_is_amo),
    .io_uop_uses_ldq(slots_12_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_12_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_12_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_12_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_12_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_12_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_12_io_uop_ldst),
    .io_uop_lrs1(slots_12_io_uop_lrs1),
    .io_uop_lrs2(slots_12_io_uop_lrs2),
    .io_uop_lrs3(slots_12_io_uop_lrs3),
    .io_uop_ldst_val(slots_12_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_12_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_12_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_12_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_12_io_uop_frs3_en),
    .io_uop_fp_val(slots_12_io_uop_fp_val),
    .io_uop_fp_single(slots_12_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_12_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_12_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_12_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_12_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_12_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_12_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_12_io_uop_debug_tsrc),
    .io_debug_p1(slots_12_io_debug_p1),
    .io_debug_p2(slots_12_io_debug_p2),
    .io_debug_p3(slots_12_io_debug_p3),
    .io_debug_ppred(slots_12_io_debug_ppred),
    .io_debug_state(slots_12_io_debug_state)
  );
  IssueSlot_16 slots_13 ( // @[issue-unit.scala 157:73]
    .clock(slots_13_clock),
    .reset(slots_13_reset),
    .io_valid(slots_13_io_valid),
    .io_will_be_valid(slots_13_io_will_be_valid),
    .io_request(slots_13_io_request),
    .io_request_hp(slots_13_io_request_hp),
    .io_grant(slots_13_io_grant),
    .io_brupdate_b1_resolve_mask(slots_13_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_13_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_13_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_13_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_13_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_13_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_13_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_13_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_13_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_13_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_13_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_13_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_13_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_13_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_13_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_13_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_13_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_13_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_13_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_13_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_13_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_13_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_13_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_13_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_13_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_13_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_13_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_13_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_13_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_13_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_13_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_13_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_13_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_13_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_13_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_13_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_13_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_13_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_13_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_13_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_13_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_13_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_13_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_13_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_13_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_13_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_13_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_13_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_13_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_13_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_13_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_13_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_13_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_13_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_13_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_13_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_13_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_13_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_13_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_13_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_13_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_13_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_13_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_13_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_13_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_13_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_13_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_13_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_13_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_13_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_13_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_13_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_13_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_13_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_13_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_13_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_13_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_13_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_13_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_13_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_13_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_13_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_13_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_13_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_13_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_13_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_13_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_13_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_13_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_13_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_13_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_13_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_13_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_13_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_13_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_13_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_13_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_13_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_13_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_13_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_13_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_13_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_13_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_13_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_13_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_13_io_brupdate_b2_target_offset),
    .io_kill(slots_13_io_kill),
    .io_clear(slots_13_io_clear),
    .io_ldspec_miss(slots_13_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_13_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_13_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_13_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_13_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_13_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_13_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_13_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_13_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_13_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_13_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_13_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_13_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_13_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_13_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_13_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_13_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_13_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_13_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_13_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_13_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_13_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_13_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_13_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_13_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_13_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_13_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_13_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_13_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_13_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_13_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_13_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_13_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_13_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_13_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_13_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_13_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_13_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_13_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_13_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_13_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_13_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_13_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_13_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_13_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_13_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_13_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_13_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_13_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_13_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_13_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_13_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_13_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_13_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_13_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_13_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_13_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_13_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_13_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_13_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_13_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_13_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_13_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_13_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_13_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_13_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_13_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_13_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_13_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_13_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_13_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_13_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_13_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_13_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_13_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_13_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_13_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_13_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_13_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_13_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_13_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_13_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_13_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_13_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_13_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_13_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_13_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_13_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_13_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_13_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_13_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_13_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_13_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_13_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_13_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_13_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_13_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_13_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_13_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_13_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_13_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_13_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_13_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_13_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_13_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_13_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_13_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_13_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_13_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_13_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_13_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_13_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_13_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_13_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_13_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_13_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_13_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_13_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_13_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_13_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_13_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_13_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_13_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_13_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_13_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_13_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_13_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_13_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_13_io_out_uop_switch),
    .io_out_uop_switch_off(slots_13_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_13_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_13_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_13_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_13_io_out_uop_rflag),
    .io_out_uop_wflag(slots_13_io_out_uop_wflag),
    .io_out_uop_prflag(slots_13_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_13_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_13_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_13_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_13_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_13_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_13_io_out_uop_split_num),
    .io_out_uop_self_index(slots_13_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_13_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_13_io_out_uop_address_num),
    .io_out_uop_uopc(slots_13_io_out_uop_uopc),
    .io_out_uop_inst(slots_13_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_13_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_13_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_13_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_13_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_13_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_13_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_13_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_13_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_13_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_13_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_13_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_13_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_13_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_13_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_13_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_13_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_13_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_13_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_13_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_13_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_13_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_13_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_13_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_13_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_13_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_13_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_13_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_13_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_13_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_13_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_13_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_13_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_13_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_13_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_13_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_13_io_out_uop_pdst),
    .io_out_uop_prs1(slots_13_io_out_uop_prs1),
    .io_out_uop_prs2(slots_13_io_out_uop_prs2),
    .io_out_uop_prs3(slots_13_io_out_uop_prs3),
    .io_out_uop_ppred(slots_13_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_13_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_13_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_13_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_13_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_13_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_13_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_13_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_13_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_13_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_13_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_13_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_13_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_13_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_13_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_13_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_13_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_13_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_13_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_13_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_13_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_13_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_13_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_13_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_13_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_13_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_13_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_13_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_13_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_13_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_13_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_13_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_13_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_13_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_13_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_13_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_13_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_13_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_13_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_13_io_uop_switch),
    .io_uop_switch_off(slots_13_io_uop_switch_off),
    .io_uop_is_unicore(slots_13_io_uop_is_unicore),
    .io_uop_shift(slots_13_io_uop_shift),
    .io_uop_lrs3_rtype(slots_13_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_13_io_uop_rflag),
    .io_uop_wflag(slots_13_io_uop_wflag),
    .io_uop_prflag(slots_13_io_uop_prflag),
    .io_uop_pwflag(slots_13_io_uop_pwflag),
    .io_uop_pflag_busy(slots_13_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_13_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_13_io_uop_op1_sel),
    .io_uop_op2_sel(slots_13_io_uop_op2_sel),
    .io_uop_split_num(slots_13_io_uop_split_num),
    .io_uop_self_index(slots_13_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_13_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_13_io_uop_address_num),
    .io_uop_uopc(slots_13_io_uop_uopc),
    .io_uop_inst(slots_13_io_uop_inst),
    .io_uop_debug_inst(slots_13_io_uop_debug_inst),
    .io_uop_is_rvc(slots_13_io_uop_is_rvc),
    .io_uop_debug_pc(slots_13_io_uop_debug_pc),
    .io_uop_iq_type(slots_13_io_uop_iq_type),
    .io_uop_fu_code(slots_13_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_13_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_13_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_13_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_13_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_13_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_13_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_13_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_13_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_13_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_13_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_13_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_13_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_13_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_13_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_13_io_uop_is_br),
    .io_uop_is_jalr(slots_13_io_uop_is_jalr),
    .io_uop_is_jal(slots_13_io_uop_is_jal),
    .io_uop_is_sfb(slots_13_io_uop_is_sfb),
    .io_uop_br_mask(slots_13_io_uop_br_mask),
    .io_uop_br_tag(slots_13_io_uop_br_tag),
    .io_uop_ftq_idx(slots_13_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_13_io_uop_edge_inst),
    .io_uop_pc_lob(slots_13_io_uop_pc_lob),
    .io_uop_taken(slots_13_io_uop_taken),
    .io_uop_imm_packed(slots_13_io_uop_imm_packed),
    .io_uop_csr_addr(slots_13_io_uop_csr_addr),
    .io_uop_rob_idx(slots_13_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_13_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_13_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_13_io_uop_rxq_idx),
    .io_uop_pdst(slots_13_io_uop_pdst),
    .io_uop_prs1(slots_13_io_uop_prs1),
    .io_uop_prs2(slots_13_io_uop_prs2),
    .io_uop_prs3(slots_13_io_uop_prs3),
    .io_uop_ppred(slots_13_io_uop_ppred),
    .io_uop_prs1_busy(slots_13_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_13_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_13_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_13_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_13_io_uop_stale_pdst),
    .io_uop_exception(slots_13_io_uop_exception),
    .io_uop_exc_cause(slots_13_io_uop_exc_cause),
    .io_uop_bypassable(slots_13_io_uop_bypassable),
    .io_uop_mem_cmd(slots_13_io_uop_mem_cmd),
    .io_uop_mem_size(slots_13_io_uop_mem_size),
    .io_uop_mem_signed(slots_13_io_uop_mem_signed),
    .io_uop_is_fence(slots_13_io_uop_is_fence),
    .io_uop_is_fencei(slots_13_io_uop_is_fencei),
    .io_uop_is_amo(slots_13_io_uop_is_amo),
    .io_uop_uses_ldq(slots_13_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_13_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_13_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_13_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_13_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_13_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_13_io_uop_ldst),
    .io_uop_lrs1(slots_13_io_uop_lrs1),
    .io_uop_lrs2(slots_13_io_uop_lrs2),
    .io_uop_lrs3(slots_13_io_uop_lrs3),
    .io_uop_ldst_val(slots_13_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_13_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_13_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_13_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_13_io_uop_frs3_en),
    .io_uop_fp_val(slots_13_io_uop_fp_val),
    .io_uop_fp_single(slots_13_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_13_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_13_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_13_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_13_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_13_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_13_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_13_io_uop_debug_tsrc),
    .io_debug_p1(slots_13_io_debug_p1),
    .io_debug_p2(slots_13_io_debug_p2),
    .io_debug_p3(slots_13_io_debug_p3),
    .io_debug_ppred(slots_13_io_debug_ppred),
    .io_debug_state(slots_13_io_debug_state)
  );
  IssueSlot_16 slots_14 ( // @[issue-unit.scala 157:73]
    .clock(slots_14_clock),
    .reset(slots_14_reset),
    .io_valid(slots_14_io_valid),
    .io_will_be_valid(slots_14_io_will_be_valid),
    .io_request(slots_14_io_request),
    .io_request_hp(slots_14_io_request_hp),
    .io_grant(slots_14_io_grant),
    .io_brupdate_b1_resolve_mask(slots_14_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_14_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_14_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_14_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_14_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_14_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_14_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_14_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_14_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_14_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_14_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_14_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_14_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_14_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_14_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_14_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_14_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_14_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_14_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_14_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_14_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_14_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_14_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_14_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_14_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_14_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_14_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_14_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_14_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_14_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_14_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_14_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_14_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_14_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_14_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_14_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_14_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_14_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_14_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_14_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_14_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_14_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_14_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_14_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_14_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_14_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_14_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_14_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_14_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_14_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_14_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_14_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_14_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_14_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_14_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_14_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_14_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_14_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_14_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_14_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_14_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_14_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_14_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_14_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_14_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_14_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_14_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_14_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_14_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_14_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_14_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_14_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_14_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_14_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_14_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_14_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_14_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_14_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_14_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_14_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_14_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_14_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_14_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_14_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_14_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_14_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_14_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_14_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_14_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_14_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_14_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_14_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_14_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_14_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_14_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_14_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_14_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_14_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_14_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_14_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_14_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_14_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_14_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_14_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_14_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_14_io_brupdate_b2_target_offset),
    .io_kill(slots_14_io_kill),
    .io_clear(slots_14_io_clear),
    .io_ldspec_miss(slots_14_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_14_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_14_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_14_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_14_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_14_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_14_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_14_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_14_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_14_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_14_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_14_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_14_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_14_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_14_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_14_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_14_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_14_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_14_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_14_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_14_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_14_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_14_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_14_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_14_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_14_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_14_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_14_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_14_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_14_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_14_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_14_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_14_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_14_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_14_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_14_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_14_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_14_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_14_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_14_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_14_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_14_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_14_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_14_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_14_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_14_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_14_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_14_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_14_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_14_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_14_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_14_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_14_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_14_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_14_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_14_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_14_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_14_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_14_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_14_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_14_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_14_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_14_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_14_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_14_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_14_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_14_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_14_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_14_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_14_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_14_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_14_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_14_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_14_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_14_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_14_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_14_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_14_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_14_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_14_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_14_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_14_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_14_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_14_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_14_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_14_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_14_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_14_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_14_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_14_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_14_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_14_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_14_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_14_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_14_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_14_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_14_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_14_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_14_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_14_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_14_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_14_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_14_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_14_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_14_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_14_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_14_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_14_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_14_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_14_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_14_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_14_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_14_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_14_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_14_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_14_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_14_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_14_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_14_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_14_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_14_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_14_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_14_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_14_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_14_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_14_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_14_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_14_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_14_io_out_uop_switch),
    .io_out_uop_switch_off(slots_14_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_14_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_14_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_14_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_14_io_out_uop_rflag),
    .io_out_uop_wflag(slots_14_io_out_uop_wflag),
    .io_out_uop_prflag(slots_14_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_14_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_14_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_14_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_14_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_14_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_14_io_out_uop_split_num),
    .io_out_uop_self_index(slots_14_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_14_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_14_io_out_uop_address_num),
    .io_out_uop_uopc(slots_14_io_out_uop_uopc),
    .io_out_uop_inst(slots_14_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_14_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_14_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_14_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_14_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_14_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_14_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_14_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_14_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_14_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_14_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_14_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_14_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_14_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_14_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_14_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_14_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_14_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_14_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_14_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_14_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_14_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_14_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_14_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_14_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_14_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_14_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_14_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_14_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_14_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_14_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_14_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_14_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_14_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_14_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_14_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_14_io_out_uop_pdst),
    .io_out_uop_prs1(slots_14_io_out_uop_prs1),
    .io_out_uop_prs2(slots_14_io_out_uop_prs2),
    .io_out_uop_prs3(slots_14_io_out_uop_prs3),
    .io_out_uop_ppred(slots_14_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_14_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_14_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_14_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_14_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_14_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_14_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_14_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_14_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_14_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_14_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_14_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_14_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_14_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_14_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_14_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_14_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_14_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_14_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_14_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_14_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_14_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_14_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_14_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_14_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_14_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_14_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_14_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_14_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_14_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_14_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_14_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_14_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_14_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_14_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_14_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_14_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_14_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_14_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_14_io_uop_switch),
    .io_uop_switch_off(slots_14_io_uop_switch_off),
    .io_uop_is_unicore(slots_14_io_uop_is_unicore),
    .io_uop_shift(slots_14_io_uop_shift),
    .io_uop_lrs3_rtype(slots_14_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_14_io_uop_rflag),
    .io_uop_wflag(slots_14_io_uop_wflag),
    .io_uop_prflag(slots_14_io_uop_prflag),
    .io_uop_pwflag(slots_14_io_uop_pwflag),
    .io_uop_pflag_busy(slots_14_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_14_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_14_io_uop_op1_sel),
    .io_uop_op2_sel(slots_14_io_uop_op2_sel),
    .io_uop_split_num(slots_14_io_uop_split_num),
    .io_uop_self_index(slots_14_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_14_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_14_io_uop_address_num),
    .io_uop_uopc(slots_14_io_uop_uopc),
    .io_uop_inst(slots_14_io_uop_inst),
    .io_uop_debug_inst(slots_14_io_uop_debug_inst),
    .io_uop_is_rvc(slots_14_io_uop_is_rvc),
    .io_uop_debug_pc(slots_14_io_uop_debug_pc),
    .io_uop_iq_type(slots_14_io_uop_iq_type),
    .io_uop_fu_code(slots_14_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_14_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_14_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_14_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_14_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_14_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_14_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_14_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_14_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_14_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_14_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_14_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_14_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_14_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_14_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_14_io_uop_is_br),
    .io_uop_is_jalr(slots_14_io_uop_is_jalr),
    .io_uop_is_jal(slots_14_io_uop_is_jal),
    .io_uop_is_sfb(slots_14_io_uop_is_sfb),
    .io_uop_br_mask(slots_14_io_uop_br_mask),
    .io_uop_br_tag(slots_14_io_uop_br_tag),
    .io_uop_ftq_idx(slots_14_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_14_io_uop_edge_inst),
    .io_uop_pc_lob(slots_14_io_uop_pc_lob),
    .io_uop_taken(slots_14_io_uop_taken),
    .io_uop_imm_packed(slots_14_io_uop_imm_packed),
    .io_uop_csr_addr(slots_14_io_uop_csr_addr),
    .io_uop_rob_idx(slots_14_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_14_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_14_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_14_io_uop_rxq_idx),
    .io_uop_pdst(slots_14_io_uop_pdst),
    .io_uop_prs1(slots_14_io_uop_prs1),
    .io_uop_prs2(slots_14_io_uop_prs2),
    .io_uop_prs3(slots_14_io_uop_prs3),
    .io_uop_ppred(slots_14_io_uop_ppred),
    .io_uop_prs1_busy(slots_14_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_14_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_14_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_14_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_14_io_uop_stale_pdst),
    .io_uop_exception(slots_14_io_uop_exception),
    .io_uop_exc_cause(slots_14_io_uop_exc_cause),
    .io_uop_bypassable(slots_14_io_uop_bypassable),
    .io_uop_mem_cmd(slots_14_io_uop_mem_cmd),
    .io_uop_mem_size(slots_14_io_uop_mem_size),
    .io_uop_mem_signed(slots_14_io_uop_mem_signed),
    .io_uop_is_fence(slots_14_io_uop_is_fence),
    .io_uop_is_fencei(slots_14_io_uop_is_fencei),
    .io_uop_is_amo(slots_14_io_uop_is_amo),
    .io_uop_uses_ldq(slots_14_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_14_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_14_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_14_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_14_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_14_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_14_io_uop_ldst),
    .io_uop_lrs1(slots_14_io_uop_lrs1),
    .io_uop_lrs2(slots_14_io_uop_lrs2),
    .io_uop_lrs3(slots_14_io_uop_lrs3),
    .io_uop_ldst_val(slots_14_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_14_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_14_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_14_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_14_io_uop_frs3_en),
    .io_uop_fp_val(slots_14_io_uop_fp_val),
    .io_uop_fp_single(slots_14_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_14_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_14_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_14_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_14_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_14_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_14_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_14_io_uop_debug_tsrc),
    .io_debug_p1(slots_14_io_debug_p1),
    .io_debug_p2(slots_14_io_debug_p2),
    .io_debug_p3(slots_14_io_debug_p3),
    .io_debug_ppred(slots_14_io_debug_ppred),
    .io_debug_state(slots_14_io_debug_state)
  );
  IssueSlot_16 slots_15 ( // @[issue-unit.scala 157:73]
    .clock(slots_15_clock),
    .reset(slots_15_reset),
    .io_valid(slots_15_io_valid),
    .io_will_be_valid(slots_15_io_will_be_valid),
    .io_request(slots_15_io_request),
    .io_request_hp(slots_15_io_request_hp),
    .io_grant(slots_15_io_grant),
    .io_brupdate_b1_resolve_mask(slots_15_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_15_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_15_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_15_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_15_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_15_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_15_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_15_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_15_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_15_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_15_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_15_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_15_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_15_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_15_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_15_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_15_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_15_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_15_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_15_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_15_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_15_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_15_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_15_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_15_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_15_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_15_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_15_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_15_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_15_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_15_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_15_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_15_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_15_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_15_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_15_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_15_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_15_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_15_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_15_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_15_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_15_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_15_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_15_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_15_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_15_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_15_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_15_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_15_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_15_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_15_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_15_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_15_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_15_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_15_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_15_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_15_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_15_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_15_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_15_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_15_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_15_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_15_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_15_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_15_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_15_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_15_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_15_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_15_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_15_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_15_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_15_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_15_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_15_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_15_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_15_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_15_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_15_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_15_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_15_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_15_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_15_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_15_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_15_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_15_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_15_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_15_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_15_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_15_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_15_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_15_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_15_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_15_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_15_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_15_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_15_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_15_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_15_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_15_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_15_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_15_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_15_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_15_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_15_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_15_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_15_io_brupdate_b2_target_offset),
    .io_kill(slots_15_io_kill),
    .io_clear(slots_15_io_clear),
    .io_ldspec_miss(slots_15_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_15_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_15_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_15_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_15_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_15_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_15_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_15_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_15_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_15_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_15_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_15_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_15_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_15_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_15_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_15_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_15_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_15_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_15_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_15_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_15_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_15_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_15_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_15_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_15_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_15_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_15_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_15_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_15_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_15_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_15_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_15_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_15_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_15_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_15_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_15_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_15_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_15_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_15_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_15_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_15_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_15_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_15_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_15_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_15_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_15_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_15_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_15_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_15_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_15_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_15_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_15_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_15_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_15_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_15_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_15_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_15_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_15_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_15_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_15_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_15_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_15_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_15_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_15_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_15_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_15_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_15_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_15_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_15_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_15_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_15_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_15_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_15_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_15_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_15_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_15_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_15_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_15_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_15_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_15_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_15_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_15_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_15_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_15_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_15_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_15_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_15_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_15_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_15_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_15_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_15_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_15_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_15_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_15_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_15_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_15_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_15_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_15_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_15_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_15_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_15_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_15_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_15_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_15_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_15_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_15_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_15_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_15_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_15_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_15_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_15_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_15_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_15_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_15_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_15_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_15_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_15_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_15_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_15_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_15_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_15_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_15_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_15_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_15_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_15_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_15_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_15_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_15_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_15_io_out_uop_switch),
    .io_out_uop_switch_off(slots_15_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_15_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_15_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_15_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_15_io_out_uop_rflag),
    .io_out_uop_wflag(slots_15_io_out_uop_wflag),
    .io_out_uop_prflag(slots_15_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_15_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_15_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_15_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_15_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_15_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_15_io_out_uop_split_num),
    .io_out_uop_self_index(slots_15_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_15_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_15_io_out_uop_address_num),
    .io_out_uop_uopc(slots_15_io_out_uop_uopc),
    .io_out_uop_inst(slots_15_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_15_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_15_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_15_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_15_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_15_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_15_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_15_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_15_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_15_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_15_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_15_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_15_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_15_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_15_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_15_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_15_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_15_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_15_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_15_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_15_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_15_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_15_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_15_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_15_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_15_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_15_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_15_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_15_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_15_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_15_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_15_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_15_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_15_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_15_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_15_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_15_io_out_uop_pdst),
    .io_out_uop_prs1(slots_15_io_out_uop_prs1),
    .io_out_uop_prs2(slots_15_io_out_uop_prs2),
    .io_out_uop_prs3(slots_15_io_out_uop_prs3),
    .io_out_uop_ppred(slots_15_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_15_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_15_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_15_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_15_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_15_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_15_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_15_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_15_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_15_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_15_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_15_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_15_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_15_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_15_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_15_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_15_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_15_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_15_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_15_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_15_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_15_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_15_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_15_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_15_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_15_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_15_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_15_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_15_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_15_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_15_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_15_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_15_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_15_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_15_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_15_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_15_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_15_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_15_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_15_io_uop_switch),
    .io_uop_switch_off(slots_15_io_uop_switch_off),
    .io_uop_is_unicore(slots_15_io_uop_is_unicore),
    .io_uop_shift(slots_15_io_uop_shift),
    .io_uop_lrs3_rtype(slots_15_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_15_io_uop_rflag),
    .io_uop_wflag(slots_15_io_uop_wflag),
    .io_uop_prflag(slots_15_io_uop_prflag),
    .io_uop_pwflag(slots_15_io_uop_pwflag),
    .io_uop_pflag_busy(slots_15_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_15_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_15_io_uop_op1_sel),
    .io_uop_op2_sel(slots_15_io_uop_op2_sel),
    .io_uop_split_num(slots_15_io_uop_split_num),
    .io_uop_self_index(slots_15_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_15_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_15_io_uop_address_num),
    .io_uop_uopc(slots_15_io_uop_uopc),
    .io_uop_inst(slots_15_io_uop_inst),
    .io_uop_debug_inst(slots_15_io_uop_debug_inst),
    .io_uop_is_rvc(slots_15_io_uop_is_rvc),
    .io_uop_debug_pc(slots_15_io_uop_debug_pc),
    .io_uop_iq_type(slots_15_io_uop_iq_type),
    .io_uop_fu_code(slots_15_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_15_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_15_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_15_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_15_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_15_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_15_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_15_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_15_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_15_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_15_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_15_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_15_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_15_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_15_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_15_io_uop_is_br),
    .io_uop_is_jalr(slots_15_io_uop_is_jalr),
    .io_uop_is_jal(slots_15_io_uop_is_jal),
    .io_uop_is_sfb(slots_15_io_uop_is_sfb),
    .io_uop_br_mask(slots_15_io_uop_br_mask),
    .io_uop_br_tag(slots_15_io_uop_br_tag),
    .io_uop_ftq_idx(slots_15_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_15_io_uop_edge_inst),
    .io_uop_pc_lob(slots_15_io_uop_pc_lob),
    .io_uop_taken(slots_15_io_uop_taken),
    .io_uop_imm_packed(slots_15_io_uop_imm_packed),
    .io_uop_csr_addr(slots_15_io_uop_csr_addr),
    .io_uop_rob_idx(slots_15_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_15_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_15_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_15_io_uop_rxq_idx),
    .io_uop_pdst(slots_15_io_uop_pdst),
    .io_uop_prs1(slots_15_io_uop_prs1),
    .io_uop_prs2(slots_15_io_uop_prs2),
    .io_uop_prs3(slots_15_io_uop_prs3),
    .io_uop_ppred(slots_15_io_uop_ppred),
    .io_uop_prs1_busy(slots_15_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_15_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_15_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_15_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_15_io_uop_stale_pdst),
    .io_uop_exception(slots_15_io_uop_exception),
    .io_uop_exc_cause(slots_15_io_uop_exc_cause),
    .io_uop_bypassable(slots_15_io_uop_bypassable),
    .io_uop_mem_cmd(slots_15_io_uop_mem_cmd),
    .io_uop_mem_size(slots_15_io_uop_mem_size),
    .io_uop_mem_signed(slots_15_io_uop_mem_signed),
    .io_uop_is_fence(slots_15_io_uop_is_fence),
    .io_uop_is_fencei(slots_15_io_uop_is_fencei),
    .io_uop_is_amo(slots_15_io_uop_is_amo),
    .io_uop_uses_ldq(slots_15_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_15_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_15_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_15_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_15_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_15_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_15_io_uop_ldst),
    .io_uop_lrs1(slots_15_io_uop_lrs1),
    .io_uop_lrs2(slots_15_io_uop_lrs2),
    .io_uop_lrs3(slots_15_io_uop_lrs3),
    .io_uop_ldst_val(slots_15_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_15_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_15_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_15_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_15_io_uop_frs3_en),
    .io_uop_fp_val(slots_15_io_uop_fp_val),
    .io_uop_fp_single(slots_15_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_15_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_15_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_15_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_15_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_15_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_15_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_15_io_uop_debug_tsrc),
    .io_debug_p1(slots_15_io_debug_p1),
    .io_debug_p2(slots_15_io_debug_p2),
    .io_debug_p3(slots_15_io_debug_p3),
    .io_debug_ppred(slots_15_io_debug_ppred),
    .io_debug_state(slots_15_io_debug_state)
  );
  IssueSlot_16 slots_16 ( // @[issue-unit.scala 157:73]
    .clock(slots_16_clock),
    .reset(slots_16_reset),
    .io_valid(slots_16_io_valid),
    .io_will_be_valid(slots_16_io_will_be_valid),
    .io_request(slots_16_io_request),
    .io_request_hp(slots_16_io_request_hp),
    .io_grant(slots_16_io_grant),
    .io_brupdate_b1_resolve_mask(slots_16_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_16_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_16_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_16_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_16_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_16_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_16_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_16_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_16_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_16_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_16_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_16_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_16_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_16_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_16_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_16_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_16_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_16_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_16_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_16_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_16_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_16_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_16_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_16_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_16_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_16_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_16_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_16_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_16_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_16_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_16_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_16_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_16_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_16_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_16_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_16_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_16_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_16_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_16_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_16_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_16_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_16_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_16_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_16_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_16_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_16_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_16_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_16_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_16_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_16_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_16_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_16_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_16_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_16_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_16_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_16_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_16_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_16_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_16_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_16_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_16_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_16_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_16_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_16_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_16_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_16_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_16_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_16_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_16_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_16_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_16_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_16_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_16_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_16_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_16_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_16_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_16_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_16_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_16_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_16_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_16_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_16_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_16_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_16_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_16_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_16_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_16_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_16_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_16_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_16_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_16_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_16_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_16_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_16_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_16_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_16_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_16_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_16_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_16_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_16_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_16_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_16_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_16_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_16_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_16_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_16_io_brupdate_b2_target_offset),
    .io_kill(slots_16_io_kill),
    .io_clear(slots_16_io_clear),
    .io_ldspec_miss(slots_16_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_16_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_16_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_16_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_16_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_16_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_16_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_16_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_16_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_16_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_16_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_16_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_16_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_16_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_16_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_16_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_16_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_16_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_16_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_16_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_16_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_16_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_16_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_16_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_16_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_16_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_16_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_16_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_16_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_16_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_16_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_16_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_16_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_16_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_16_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_16_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_16_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_16_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_16_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_16_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_16_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_16_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_16_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_16_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_16_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_16_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_16_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_16_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_16_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_16_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_16_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_16_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_16_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_16_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_16_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_16_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_16_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_16_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_16_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_16_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_16_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_16_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_16_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_16_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_16_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_16_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_16_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_16_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_16_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_16_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_16_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_16_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_16_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_16_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_16_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_16_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_16_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_16_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_16_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_16_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_16_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_16_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_16_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_16_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_16_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_16_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_16_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_16_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_16_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_16_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_16_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_16_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_16_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_16_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_16_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_16_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_16_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_16_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_16_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_16_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_16_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_16_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_16_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_16_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_16_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_16_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_16_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_16_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_16_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_16_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_16_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_16_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_16_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_16_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_16_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_16_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_16_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_16_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_16_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_16_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_16_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_16_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_16_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_16_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_16_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_16_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_16_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_16_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_16_io_out_uop_switch),
    .io_out_uop_switch_off(slots_16_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_16_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_16_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_16_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_16_io_out_uop_rflag),
    .io_out_uop_wflag(slots_16_io_out_uop_wflag),
    .io_out_uop_prflag(slots_16_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_16_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_16_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_16_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_16_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_16_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_16_io_out_uop_split_num),
    .io_out_uop_self_index(slots_16_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_16_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_16_io_out_uop_address_num),
    .io_out_uop_uopc(slots_16_io_out_uop_uopc),
    .io_out_uop_inst(slots_16_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_16_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_16_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_16_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_16_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_16_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_16_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_16_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_16_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_16_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_16_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_16_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_16_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_16_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_16_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_16_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_16_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_16_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_16_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_16_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_16_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_16_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_16_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_16_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_16_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_16_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_16_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_16_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_16_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_16_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_16_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_16_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_16_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_16_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_16_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_16_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_16_io_out_uop_pdst),
    .io_out_uop_prs1(slots_16_io_out_uop_prs1),
    .io_out_uop_prs2(slots_16_io_out_uop_prs2),
    .io_out_uop_prs3(slots_16_io_out_uop_prs3),
    .io_out_uop_ppred(slots_16_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_16_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_16_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_16_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_16_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_16_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_16_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_16_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_16_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_16_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_16_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_16_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_16_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_16_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_16_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_16_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_16_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_16_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_16_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_16_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_16_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_16_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_16_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_16_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_16_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_16_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_16_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_16_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_16_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_16_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_16_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_16_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_16_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_16_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_16_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_16_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_16_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_16_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_16_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_16_io_uop_switch),
    .io_uop_switch_off(slots_16_io_uop_switch_off),
    .io_uop_is_unicore(slots_16_io_uop_is_unicore),
    .io_uop_shift(slots_16_io_uop_shift),
    .io_uop_lrs3_rtype(slots_16_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_16_io_uop_rflag),
    .io_uop_wflag(slots_16_io_uop_wflag),
    .io_uop_prflag(slots_16_io_uop_prflag),
    .io_uop_pwflag(slots_16_io_uop_pwflag),
    .io_uop_pflag_busy(slots_16_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_16_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_16_io_uop_op1_sel),
    .io_uop_op2_sel(slots_16_io_uop_op2_sel),
    .io_uop_split_num(slots_16_io_uop_split_num),
    .io_uop_self_index(slots_16_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_16_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_16_io_uop_address_num),
    .io_uop_uopc(slots_16_io_uop_uopc),
    .io_uop_inst(slots_16_io_uop_inst),
    .io_uop_debug_inst(slots_16_io_uop_debug_inst),
    .io_uop_is_rvc(slots_16_io_uop_is_rvc),
    .io_uop_debug_pc(slots_16_io_uop_debug_pc),
    .io_uop_iq_type(slots_16_io_uop_iq_type),
    .io_uop_fu_code(slots_16_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_16_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_16_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_16_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_16_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_16_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_16_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_16_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_16_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_16_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_16_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_16_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_16_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_16_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_16_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_16_io_uop_is_br),
    .io_uop_is_jalr(slots_16_io_uop_is_jalr),
    .io_uop_is_jal(slots_16_io_uop_is_jal),
    .io_uop_is_sfb(slots_16_io_uop_is_sfb),
    .io_uop_br_mask(slots_16_io_uop_br_mask),
    .io_uop_br_tag(slots_16_io_uop_br_tag),
    .io_uop_ftq_idx(slots_16_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_16_io_uop_edge_inst),
    .io_uop_pc_lob(slots_16_io_uop_pc_lob),
    .io_uop_taken(slots_16_io_uop_taken),
    .io_uop_imm_packed(slots_16_io_uop_imm_packed),
    .io_uop_csr_addr(slots_16_io_uop_csr_addr),
    .io_uop_rob_idx(slots_16_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_16_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_16_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_16_io_uop_rxq_idx),
    .io_uop_pdst(slots_16_io_uop_pdst),
    .io_uop_prs1(slots_16_io_uop_prs1),
    .io_uop_prs2(slots_16_io_uop_prs2),
    .io_uop_prs3(slots_16_io_uop_prs3),
    .io_uop_ppred(slots_16_io_uop_ppred),
    .io_uop_prs1_busy(slots_16_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_16_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_16_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_16_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_16_io_uop_stale_pdst),
    .io_uop_exception(slots_16_io_uop_exception),
    .io_uop_exc_cause(slots_16_io_uop_exc_cause),
    .io_uop_bypassable(slots_16_io_uop_bypassable),
    .io_uop_mem_cmd(slots_16_io_uop_mem_cmd),
    .io_uop_mem_size(slots_16_io_uop_mem_size),
    .io_uop_mem_signed(slots_16_io_uop_mem_signed),
    .io_uop_is_fence(slots_16_io_uop_is_fence),
    .io_uop_is_fencei(slots_16_io_uop_is_fencei),
    .io_uop_is_amo(slots_16_io_uop_is_amo),
    .io_uop_uses_ldq(slots_16_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_16_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_16_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_16_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_16_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_16_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_16_io_uop_ldst),
    .io_uop_lrs1(slots_16_io_uop_lrs1),
    .io_uop_lrs2(slots_16_io_uop_lrs2),
    .io_uop_lrs3(slots_16_io_uop_lrs3),
    .io_uop_ldst_val(slots_16_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_16_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_16_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_16_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_16_io_uop_frs3_en),
    .io_uop_fp_val(slots_16_io_uop_fp_val),
    .io_uop_fp_single(slots_16_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_16_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_16_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_16_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_16_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_16_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_16_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_16_io_uop_debug_tsrc),
    .io_debug_p1(slots_16_io_debug_p1),
    .io_debug_p2(slots_16_io_debug_p2),
    .io_debug_p3(slots_16_io_debug_p3),
    .io_debug_ppred(slots_16_io_debug_ppred),
    .io_debug_state(slots_16_io_debug_state)
  );
  IssueSlot_16 slots_17 ( // @[issue-unit.scala 157:73]
    .clock(slots_17_clock),
    .reset(slots_17_reset),
    .io_valid(slots_17_io_valid),
    .io_will_be_valid(slots_17_io_will_be_valid),
    .io_request(slots_17_io_request),
    .io_request_hp(slots_17_io_request_hp),
    .io_grant(slots_17_io_grant),
    .io_brupdate_b1_resolve_mask(slots_17_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_17_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_17_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_17_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_17_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_17_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_17_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_17_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_17_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_17_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_17_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_17_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_17_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_17_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_17_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_17_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_17_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_17_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_17_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_17_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_17_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_17_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_17_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_17_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_17_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_17_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_17_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_17_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_17_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_17_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_17_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_17_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_17_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_17_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_17_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_17_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_17_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_17_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_17_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_17_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_17_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_17_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_17_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_17_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_17_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_17_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_17_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_17_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_17_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_17_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_17_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_17_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_17_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_17_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_17_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_17_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_17_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_17_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_17_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_17_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_17_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_17_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_17_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_17_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_17_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_17_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_17_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_17_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_17_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_17_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_17_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_17_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_17_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_17_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_17_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_17_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_17_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_17_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_17_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_17_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_17_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_17_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_17_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_17_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_17_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_17_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_17_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_17_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_17_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_17_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_17_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_17_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_17_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_17_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_17_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_17_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_17_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_17_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_17_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_17_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_17_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_17_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_17_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_17_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_17_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_17_io_brupdate_b2_target_offset),
    .io_kill(slots_17_io_kill),
    .io_clear(slots_17_io_clear),
    .io_ldspec_miss(slots_17_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_17_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_17_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_17_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_17_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_17_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_17_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_17_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_17_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_17_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_17_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_17_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_17_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_17_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_17_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_17_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_17_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_17_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_17_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_17_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_17_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_17_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_17_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_17_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_17_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_17_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_17_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_17_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_17_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_17_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_17_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_17_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_17_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_17_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_17_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_17_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_17_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_17_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_17_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_17_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_17_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_17_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_17_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_17_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_17_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_17_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_17_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_17_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_17_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_17_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_17_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_17_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_17_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_17_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_17_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_17_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_17_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_17_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_17_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_17_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_17_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_17_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_17_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_17_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_17_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_17_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_17_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_17_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_17_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_17_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_17_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_17_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_17_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_17_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_17_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_17_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_17_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_17_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_17_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_17_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_17_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_17_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_17_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_17_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_17_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_17_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_17_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_17_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_17_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_17_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_17_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_17_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_17_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_17_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_17_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_17_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_17_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_17_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_17_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_17_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_17_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_17_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_17_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_17_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_17_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_17_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_17_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_17_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_17_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_17_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_17_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_17_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_17_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_17_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_17_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_17_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_17_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_17_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_17_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_17_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_17_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_17_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_17_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_17_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_17_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_17_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_17_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_17_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_17_io_out_uop_switch),
    .io_out_uop_switch_off(slots_17_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_17_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_17_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_17_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_17_io_out_uop_rflag),
    .io_out_uop_wflag(slots_17_io_out_uop_wflag),
    .io_out_uop_prflag(slots_17_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_17_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_17_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_17_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_17_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_17_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_17_io_out_uop_split_num),
    .io_out_uop_self_index(slots_17_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_17_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_17_io_out_uop_address_num),
    .io_out_uop_uopc(slots_17_io_out_uop_uopc),
    .io_out_uop_inst(slots_17_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_17_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_17_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_17_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_17_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_17_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_17_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_17_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_17_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_17_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_17_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_17_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_17_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_17_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_17_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_17_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_17_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_17_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_17_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_17_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_17_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_17_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_17_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_17_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_17_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_17_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_17_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_17_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_17_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_17_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_17_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_17_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_17_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_17_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_17_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_17_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_17_io_out_uop_pdst),
    .io_out_uop_prs1(slots_17_io_out_uop_prs1),
    .io_out_uop_prs2(slots_17_io_out_uop_prs2),
    .io_out_uop_prs3(slots_17_io_out_uop_prs3),
    .io_out_uop_ppred(slots_17_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_17_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_17_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_17_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_17_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_17_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_17_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_17_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_17_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_17_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_17_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_17_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_17_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_17_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_17_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_17_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_17_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_17_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_17_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_17_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_17_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_17_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_17_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_17_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_17_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_17_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_17_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_17_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_17_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_17_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_17_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_17_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_17_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_17_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_17_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_17_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_17_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_17_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_17_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_17_io_uop_switch),
    .io_uop_switch_off(slots_17_io_uop_switch_off),
    .io_uop_is_unicore(slots_17_io_uop_is_unicore),
    .io_uop_shift(slots_17_io_uop_shift),
    .io_uop_lrs3_rtype(slots_17_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_17_io_uop_rflag),
    .io_uop_wflag(slots_17_io_uop_wflag),
    .io_uop_prflag(slots_17_io_uop_prflag),
    .io_uop_pwflag(slots_17_io_uop_pwflag),
    .io_uop_pflag_busy(slots_17_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_17_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_17_io_uop_op1_sel),
    .io_uop_op2_sel(slots_17_io_uop_op2_sel),
    .io_uop_split_num(slots_17_io_uop_split_num),
    .io_uop_self_index(slots_17_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_17_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_17_io_uop_address_num),
    .io_uop_uopc(slots_17_io_uop_uopc),
    .io_uop_inst(slots_17_io_uop_inst),
    .io_uop_debug_inst(slots_17_io_uop_debug_inst),
    .io_uop_is_rvc(slots_17_io_uop_is_rvc),
    .io_uop_debug_pc(slots_17_io_uop_debug_pc),
    .io_uop_iq_type(slots_17_io_uop_iq_type),
    .io_uop_fu_code(slots_17_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_17_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_17_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_17_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_17_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_17_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_17_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_17_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_17_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_17_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_17_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_17_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_17_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_17_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_17_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_17_io_uop_is_br),
    .io_uop_is_jalr(slots_17_io_uop_is_jalr),
    .io_uop_is_jal(slots_17_io_uop_is_jal),
    .io_uop_is_sfb(slots_17_io_uop_is_sfb),
    .io_uop_br_mask(slots_17_io_uop_br_mask),
    .io_uop_br_tag(slots_17_io_uop_br_tag),
    .io_uop_ftq_idx(slots_17_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_17_io_uop_edge_inst),
    .io_uop_pc_lob(slots_17_io_uop_pc_lob),
    .io_uop_taken(slots_17_io_uop_taken),
    .io_uop_imm_packed(slots_17_io_uop_imm_packed),
    .io_uop_csr_addr(slots_17_io_uop_csr_addr),
    .io_uop_rob_idx(slots_17_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_17_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_17_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_17_io_uop_rxq_idx),
    .io_uop_pdst(slots_17_io_uop_pdst),
    .io_uop_prs1(slots_17_io_uop_prs1),
    .io_uop_prs2(slots_17_io_uop_prs2),
    .io_uop_prs3(slots_17_io_uop_prs3),
    .io_uop_ppred(slots_17_io_uop_ppred),
    .io_uop_prs1_busy(slots_17_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_17_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_17_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_17_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_17_io_uop_stale_pdst),
    .io_uop_exception(slots_17_io_uop_exception),
    .io_uop_exc_cause(slots_17_io_uop_exc_cause),
    .io_uop_bypassable(slots_17_io_uop_bypassable),
    .io_uop_mem_cmd(slots_17_io_uop_mem_cmd),
    .io_uop_mem_size(slots_17_io_uop_mem_size),
    .io_uop_mem_signed(slots_17_io_uop_mem_signed),
    .io_uop_is_fence(slots_17_io_uop_is_fence),
    .io_uop_is_fencei(slots_17_io_uop_is_fencei),
    .io_uop_is_amo(slots_17_io_uop_is_amo),
    .io_uop_uses_ldq(slots_17_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_17_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_17_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_17_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_17_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_17_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_17_io_uop_ldst),
    .io_uop_lrs1(slots_17_io_uop_lrs1),
    .io_uop_lrs2(slots_17_io_uop_lrs2),
    .io_uop_lrs3(slots_17_io_uop_lrs3),
    .io_uop_ldst_val(slots_17_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_17_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_17_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_17_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_17_io_uop_frs3_en),
    .io_uop_fp_val(slots_17_io_uop_fp_val),
    .io_uop_fp_single(slots_17_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_17_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_17_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_17_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_17_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_17_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_17_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_17_io_uop_debug_tsrc),
    .io_debug_p1(slots_17_io_debug_p1),
    .io_debug_p2(slots_17_io_debug_p2),
    .io_debug_p3(slots_17_io_debug_p3),
    .io_debug_ppred(slots_17_io_debug_ppred),
    .io_debug_state(slots_17_io_debug_state)
  );
  IssueSlot_16 slots_18 ( // @[issue-unit.scala 157:73]
    .clock(slots_18_clock),
    .reset(slots_18_reset),
    .io_valid(slots_18_io_valid),
    .io_will_be_valid(slots_18_io_will_be_valid),
    .io_request(slots_18_io_request),
    .io_request_hp(slots_18_io_request_hp),
    .io_grant(slots_18_io_grant),
    .io_brupdate_b1_resolve_mask(slots_18_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_18_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_18_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_18_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_18_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_18_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_18_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_18_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_18_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_18_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_18_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_18_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_18_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_18_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_18_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_18_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_18_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_18_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_18_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_18_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_18_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_18_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_18_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_18_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_18_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_18_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_18_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_18_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_18_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_18_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_18_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_18_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_18_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_18_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_18_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_18_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_18_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_18_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_18_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_18_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_18_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_18_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_18_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_18_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_18_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_18_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_18_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_18_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_18_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_18_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_18_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_18_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_18_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_18_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_18_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_18_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_18_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_18_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_18_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_18_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_18_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_18_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_18_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_18_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_18_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_18_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_18_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_18_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_18_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_18_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_18_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_18_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_18_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_18_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_18_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_18_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_18_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_18_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_18_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_18_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_18_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_18_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_18_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_18_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_18_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_18_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_18_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_18_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_18_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_18_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_18_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_18_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_18_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_18_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_18_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_18_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_18_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_18_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_18_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_18_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_18_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_18_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_18_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_18_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_18_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_18_io_brupdate_b2_target_offset),
    .io_kill(slots_18_io_kill),
    .io_clear(slots_18_io_clear),
    .io_ldspec_miss(slots_18_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_18_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_18_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_18_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_18_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_18_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_18_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_18_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_18_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_18_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_18_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_18_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_18_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_18_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_18_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_18_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_18_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_18_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_18_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_18_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_18_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_18_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_18_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_18_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_18_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_18_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_18_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_18_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_18_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_18_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_18_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_18_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_18_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_18_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_18_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_18_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_18_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_18_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_18_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_18_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_18_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_18_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_18_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_18_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_18_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_18_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_18_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_18_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_18_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_18_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_18_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_18_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_18_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_18_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_18_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_18_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_18_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_18_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_18_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_18_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_18_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_18_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_18_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_18_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_18_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_18_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_18_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_18_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_18_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_18_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_18_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_18_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_18_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_18_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_18_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_18_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_18_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_18_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_18_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_18_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_18_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_18_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_18_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_18_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_18_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_18_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_18_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_18_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_18_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_18_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_18_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_18_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_18_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_18_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_18_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_18_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_18_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_18_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_18_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_18_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_18_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_18_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_18_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_18_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_18_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_18_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_18_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_18_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_18_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_18_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_18_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_18_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_18_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_18_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_18_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_18_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_18_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_18_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_18_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_18_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_18_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_18_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_18_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_18_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_18_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_18_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_18_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_18_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_18_io_out_uop_switch),
    .io_out_uop_switch_off(slots_18_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_18_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_18_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_18_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_18_io_out_uop_rflag),
    .io_out_uop_wflag(slots_18_io_out_uop_wflag),
    .io_out_uop_prflag(slots_18_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_18_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_18_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_18_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_18_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_18_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_18_io_out_uop_split_num),
    .io_out_uop_self_index(slots_18_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_18_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_18_io_out_uop_address_num),
    .io_out_uop_uopc(slots_18_io_out_uop_uopc),
    .io_out_uop_inst(slots_18_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_18_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_18_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_18_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_18_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_18_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_18_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_18_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_18_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_18_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_18_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_18_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_18_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_18_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_18_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_18_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_18_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_18_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_18_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_18_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_18_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_18_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_18_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_18_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_18_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_18_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_18_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_18_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_18_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_18_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_18_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_18_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_18_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_18_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_18_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_18_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_18_io_out_uop_pdst),
    .io_out_uop_prs1(slots_18_io_out_uop_prs1),
    .io_out_uop_prs2(slots_18_io_out_uop_prs2),
    .io_out_uop_prs3(slots_18_io_out_uop_prs3),
    .io_out_uop_ppred(slots_18_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_18_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_18_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_18_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_18_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_18_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_18_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_18_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_18_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_18_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_18_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_18_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_18_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_18_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_18_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_18_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_18_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_18_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_18_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_18_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_18_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_18_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_18_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_18_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_18_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_18_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_18_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_18_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_18_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_18_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_18_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_18_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_18_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_18_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_18_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_18_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_18_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_18_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_18_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_18_io_uop_switch),
    .io_uop_switch_off(slots_18_io_uop_switch_off),
    .io_uop_is_unicore(slots_18_io_uop_is_unicore),
    .io_uop_shift(slots_18_io_uop_shift),
    .io_uop_lrs3_rtype(slots_18_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_18_io_uop_rflag),
    .io_uop_wflag(slots_18_io_uop_wflag),
    .io_uop_prflag(slots_18_io_uop_prflag),
    .io_uop_pwflag(slots_18_io_uop_pwflag),
    .io_uop_pflag_busy(slots_18_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_18_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_18_io_uop_op1_sel),
    .io_uop_op2_sel(slots_18_io_uop_op2_sel),
    .io_uop_split_num(slots_18_io_uop_split_num),
    .io_uop_self_index(slots_18_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_18_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_18_io_uop_address_num),
    .io_uop_uopc(slots_18_io_uop_uopc),
    .io_uop_inst(slots_18_io_uop_inst),
    .io_uop_debug_inst(slots_18_io_uop_debug_inst),
    .io_uop_is_rvc(slots_18_io_uop_is_rvc),
    .io_uop_debug_pc(slots_18_io_uop_debug_pc),
    .io_uop_iq_type(slots_18_io_uop_iq_type),
    .io_uop_fu_code(slots_18_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_18_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_18_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_18_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_18_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_18_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_18_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_18_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_18_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_18_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_18_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_18_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_18_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_18_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_18_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_18_io_uop_is_br),
    .io_uop_is_jalr(slots_18_io_uop_is_jalr),
    .io_uop_is_jal(slots_18_io_uop_is_jal),
    .io_uop_is_sfb(slots_18_io_uop_is_sfb),
    .io_uop_br_mask(slots_18_io_uop_br_mask),
    .io_uop_br_tag(slots_18_io_uop_br_tag),
    .io_uop_ftq_idx(slots_18_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_18_io_uop_edge_inst),
    .io_uop_pc_lob(slots_18_io_uop_pc_lob),
    .io_uop_taken(slots_18_io_uop_taken),
    .io_uop_imm_packed(slots_18_io_uop_imm_packed),
    .io_uop_csr_addr(slots_18_io_uop_csr_addr),
    .io_uop_rob_idx(slots_18_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_18_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_18_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_18_io_uop_rxq_idx),
    .io_uop_pdst(slots_18_io_uop_pdst),
    .io_uop_prs1(slots_18_io_uop_prs1),
    .io_uop_prs2(slots_18_io_uop_prs2),
    .io_uop_prs3(slots_18_io_uop_prs3),
    .io_uop_ppred(slots_18_io_uop_ppred),
    .io_uop_prs1_busy(slots_18_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_18_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_18_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_18_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_18_io_uop_stale_pdst),
    .io_uop_exception(slots_18_io_uop_exception),
    .io_uop_exc_cause(slots_18_io_uop_exc_cause),
    .io_uop_bypassable(slots_18_io_uop_bypassable),
    .io_uop_mem_cmd(slots_18_io_uop_mem_cmd),
    .io_uop_mem_size(slots_18_io_uop_mem_size),
    .io_uop_mem_signed(slots_18_io_uop_mem_signed),
    .io_uop_is_fence(slots_18_io_uop_is_fence),
    .io_uop_is_fencei(slots_18_io_uop_is_fencei),
    .io_uop_is_amo(slots_18_io_uop_is_amo),
    .io_uop_uses_ldq(slots_18_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_18_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_18_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_18_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_18_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_18_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_18_io_uop_ldst),
    .io_uop_lrs1(slots_18_io_uop_lrs1),
    .io_uop_lrs2(slots_18_io_uop_lrs2),
    .io_uop_lrs3(slots_18_io_uop_lrs3),
    .io_uop_ldst_val(slots_18_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_18_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_18_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_18_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_18_io_uop_frs3_en),
    .io_uop_fp_val(slots_18_io_uop_fp_val),
    .io_uop_fp_single(slots_18_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_18_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_18_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_18_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_18_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_18_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_18_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_18_io_uop_debug_tsrc),
    .io_debug_p1(slots_18_io_debug_p1),
    .io_debug_p2(slots_18_io_debug_p2),
    .io_debug_p3(slots_18_io_debug_p3),
    .io_debug_ppred(slots_18_io_debug_ppred),
    .io_debug_state(slots_18_io_debug_state)
  );
  IssueSlot_16 slots_19 ( // @[issue-unit.scala 157:73]
    .clock(slots_19_clock),
    .reset(slots_19_reset),
    .io_valid(slots_19_io_valid),
    .io_will_be_valid(slots_19_io_will_be_valid),
    .io_request(slots_19_io_request),
    .io_request_hp(slots_19_io_request_hp),
    .io_grant(slots_19_io_grant),
    .io_brupdate_b1_resolve_mask(slots_19_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_19_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_19_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_19_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_19_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_19_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_19_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_19_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_19_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_19_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_19_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_19_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_19_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_19_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_19_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_19_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_19_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_19_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_19_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_19_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_19_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_19_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_19_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_19_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_19_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_19_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_19_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_19_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_19_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_19_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_19_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_19_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_19_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_19_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_19_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_19_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_19_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_19_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_19_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_19_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_19_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_19_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_19_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_19_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_19_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_19_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_19_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_19_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_19_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_19_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_19_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_19_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_19_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_19_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_19_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_19_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_19_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_19_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_19_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_19_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_19_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_19_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_19_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_19_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_19_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_19_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_19_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_19_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_19_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_19_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_19_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_19_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_19_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_19_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_19_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_19_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_19_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_19_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_19_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_19_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_19_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_19_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_19_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_19_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_19_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_19_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_19_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_19_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_19_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_19_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_19_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_19_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_19_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_19_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_19_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_19_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_19_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_19_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_19_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_19_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_19_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_19_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_19_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_19_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_19_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_19_io_brupdate_b2_target_offset),
    .io_kill(slots_19_io_kill),
    .io_clear(slots_19_io_clear),
    .io_ldspec_miss(slots_19_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_19_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_19_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_19_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_19_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_19_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_19_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_19_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_19_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_19_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_19_io_wakeup_ports_1_bits_flag_valid),
    .io_wakeup_ports_2_valid(slots_19_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_19_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_19_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_2_bits_pwflag(slots_19_io_wakeup_ports_2_bits_pwflag),
    .io_wakeup_ports_2_bits_flag_valid(slots_19_io_wakeup_ports_2_bits_flag_valid),
    .io_wakeup_ports_3_valid(slots_19_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_19_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_19_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_3_bits_pwflag(slots_19_io_wakeup_ports_3_bits_pwflag),
    .io_wakeup_ports_3_bits_flag_valid(slots_19_io_wakeup_ports_3_bits_flag_valid),
    .io_wakeup_ports_4_valid(slots_19_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_19_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_19_io_wakeup_ports_4_bits_poisoned),
    .io_wakeup_ports_4_bits_pwflag(slots_19_io_wakeup_ports_4_bits_pwflag),
    .io_wakeup_ports_4_bits_flag_valid(slots_19_io_wakeup_ports_4_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_19_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_19_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_19_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_19_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_19_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_19_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_19_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_19_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_19_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_19_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_19_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_19_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_19_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_19_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_19_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_19_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_19_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_19_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_19_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_19_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_19_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_19_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_19_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_19_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_19_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_19_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_19_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_19_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_19_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_19_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_19_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_19_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_19_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_19_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_19_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_19_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_19_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_19_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_19_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_19_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_19_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_19_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_19_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_19_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_19_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_19_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_19_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_19_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_19_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_19_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_19_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_19_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_19_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_19_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_19_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_19_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_19_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_19_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_19_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_19_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_19_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_19_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_19_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_19_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_19_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_19_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_19_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_19_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_19_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_19_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_19_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_19_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_19_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_19_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_19_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_19_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_19_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_19_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_19_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_19_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_19_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_19_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_19_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_19_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_19_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_19_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_19_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_19_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_19_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_19_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_19_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_19_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_19_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_19_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_19_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_19_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_19_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_19_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_19_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_19_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_19_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_19_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_19_io_out_uop_switch),
    .io_out_uop_switch_off(slots_19_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_19_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_19_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_19_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_19_io_out_uop_rflag),
    .io_out_uop_wflag(slots_19_io_out_uop_wflag),
    .io_out_uop_prflag(slots_19_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_19_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_19_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_19_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_19_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_19_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_19_io_out_uop_split_num),
    .io_out_uop_self_index(slots_19_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_19_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_19_io_out_uop_address_num),
    .io_out_uop_uopc(slots_19_io_out_uop_uopc),
    .io_out_uop_inst(slots_19_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_19_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_19_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_19_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_19_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_19_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_19_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_19_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_19_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_19_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_19_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_19_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_19_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_19_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_19_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_19_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_19_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_19_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_19_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_19_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_19_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_19_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_19_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_19_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_19_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_19_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_19_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_19_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_19_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_19_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_19_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_19_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_19_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_19_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_19_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_19_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_19_io_out_uop_pdst),
    .io_out_uop_prs1(slots_19_io_out_uop_prs1),
    .io_out_uop_prs2(slots_19_io_out_uop_prs2),
    .io_out_uop_prs3(slots_19_io_out_uop_prs3),
    .io_out_uop_ppred(slots_19_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_19_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_19_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_19_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_19_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_19_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_19_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_19_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_19_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_19_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_19_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_19_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_19_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_19_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_19_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_19_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_19_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_19_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_19_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_19_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_19_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_19_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_19_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_19_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_19_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_19_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_19_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_19_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_19_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_19_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_19_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_19_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_19_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_19_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_19_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_19_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_19_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_19_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_19_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_19_io_uop_switch),
    .io_uop_switch_off(slots_19_io_uop_switch_off),
    .io_uop_is_unicore(slots_19_io_uop_is_unicore),
    .io_uop_shift(slots_19_io_uop_shift),
    .io_uop_lrs3_rtype(slots_19_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_19_io_uop_rflag),
    .io_uop_wflag(slots_19_io_uop_wflag),
    .io_uop_prflag(slots_19_io_uop_prflag),
    .io_uop_pwflag(slots_19_io_uop_pwflag),
    .io_uop_pflag_busy(slots_19_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_19_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_19_io_uop_op1_sel),
    .io_uop_op2_sel(slots_19_io_uop_op2_sel),
    .io_uop_split_num(slots_19_io_uop_split_num),
    .io_uop_self_index(slots_19_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_19_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_19_io_uop_address_num),
    .io_uop_uopc(slots_19_io_uop_uopc),
    .io_uop_inst(slots_19_io_uop_inst),
    .io_uop_debug_inst(slots_19_io_uop_debug_inst),
    .io_uop_is_rvc(slots_19_io_uop_is_rvc),
    .io_uop_debug_pc(slots_19_io_uop_debug_pc),
    .io_uop_iq_type(slots_19_io_uop_iq_type),
    .io_uop_fu_code(slots_19_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_19_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_19_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_19_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_19_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_19_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_19_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_19_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_19_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_19_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_19_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_19_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_19_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_19_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_19_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_19_io_uop_is_br),
    .io_uop_is_jalr(slots_19_io_uop_is_jalr),
    .io_uop_is_jal(slots_19_io_uop_is_jal),
    .io_uop_is_sfb(slots_19_io_uop_is_sfb),
    .io_uop_br_mask(slots_19_io_uop_br_mask),
    .io_uop_br_tag(slots_19_io_uop_br_tag),
    .io_uop_ftq_idx(slots_19_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_19_io_uop_edge_inst),
    .io_uop_pc_lob(slots_19_io_uop_pc_lob),
    .io_uop_taken(slots_19_io_uop_taken),
    .io_uop_imm_packed(slots_19_io_uop_imm_packed),
    .io_uop_csr_addr(slots_19_io_uop_csr_addr),
    .io_uop_rob_idx(slots_19_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_19_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_19_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_19_io_uop_rxq_idx),
    .io_uop_pdst(slots_19_io_uop_pdst),
    .io_uop_prs1(slots_19_io_uop_prs1),
    .io_uop_prs2(slots_19_io_uop_prs2),
    .io_uop_prs3(slots_19_io_uop_prs3),
    .io_uop_ppred(slots_19_io_uop_ppred),
    .io_uop_prs1_busy(slots_19_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_19_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_19_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_19_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_19_io_uop_stale_pdst),
    .io_uop_exception(slots_19_io_uop_exception),
    .io_uop_exc_cause(slots_19_io_uop_exc_cause),
    .io_uop_bypassable(slots_19_io_uop_bypassable),
    .io_uop_mem_cmd(slots_19_io_uop_mem_cmd),
    .io_uop_mem_size(slots_19_io_uop_mem_size),
    .io_uop_mem_signed(slots_19_io_uop_mem_signed),
    .io_uop_is_fence(slots_19_io_uop_is_fence),
    .io_uop_is_fencei(slots_19_io_uop_is_fencei),
    .io_uop_is_amo(slots_19_io_uop_is_amo),
    .io_uop_uses_ldq(slots_19_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_19_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_19_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_19_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_19_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_19_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_19_io_uop_ldst),
    .io_uop_lrs1(slots_19_io_uop_lrs1),
    .io_uop_lrs2(slots_19_io_uop_lrs2),
    .io_uop_lrs3(slots_19_io_uop_lrs3),
    .io_uop_ldst_val(slots_19_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_19_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_19_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_19_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_19_io_uop_frs3_en),
    .io_uop_fp_val(slots_19_io_uop_fp_val),
    .io_uop_fp_single(slots_19_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_19_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_19_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_19_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_19_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_19_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_19_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_19_io_uop_debug_tsrc),
    .io_debug_p1(slots_19_io_debug_p1),
    .io_debug_p2(slots_19_io_debug_p2),
    .io_debug_p3(slots_19_io_debug_p3),
    .io_debug_ppred(slots_19_io_debug_ppred),
    .io_debug_state(slots_19_io_debug_state)
  );
  assign io_dis_uops_0_ready = REG; // @[issue-unit-age-ordered.scala 87:26]
  assign io_dis_uops_1_ready = REG_1; // @[issue-unit-age-ordered.scala 87:26]
  assign io_iss_valids_0 = _T_995 | (_T_965 | (_T_935 | (_T_905 | (_T_875 | (_T_845 | (_T_815 | (_T_785 | (_T_755 | (
    _T_725 | (_T_695 | (_T_665 | (_T_635 | (_T_605 | (_T_575 | (_T_545 | (_T_515 | (_T_485 | (_T_455 | _T_423)))))))))))
    ))))))); // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 124:26]
  assign io_iss_valids_1 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 | (issue_slots_18_request & ~_T_965 &
    _T_968 & ~_T_947 | (_T_946 & ~_T_917 | (issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 | (
    issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 | _GEN_6843)))); // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 124:26]
  assign io_iss_uops_0_switch = _T_995 ? issue_slots_19_uop_switch : _GEN_7633; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_switch_off = _T_995 ? issue_slots_19_uop_switch_off : _GEN_7632; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_unicore = _T_995 ? issue_slots_19_uop_is_unicore : _GEN_7631; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_shift = _T_995 ? issue_slots_19_uop_shift : _GEN_7630; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs3_rtype = _T_995 ? issue_slots_19_uop_lrs3_rtype : _GEN_7629; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rflag = _T_995 ? issue_slots_19_uop_rflag : _GEN_7628; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_wflag = _T_995 ? issue_slots_19_uop_wflag : _GEN_7627; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prflag = _T_995 ? issue_slots_19_uop_prflag : _GEN_7626; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pwflag = _T_995 ? issue_slots_19_uop_pwflag : _GEN_7625; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pflag_busy = _T_995 ? issue_slots_19_uop_pflag_busy : _GEN_7624; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_stale_pflag = _T_995 ? issue_slots_19_uop_stale_pflag : _GEN_7623; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_op1_sel = _T_995 ? issue_slots_19_uop_op1_sel : _GEN_7622; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_op2_sel = _T_995 ? issue_slots_19_uop_op2_sel : _GEN_7621; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_split_num = _T_995 ? issue_slots_19_uop_split_num : _GEN_7620; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_self_index = _T_995 ? issue_slots_19_uop_self_index : _GEN_7619; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rob_inst_idx = _T_995 ? issue_slots_19_uop_rob_inst_idx : _GEN_7618; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_address_num = _T_995 ? issue_slots_19_uop_address_num : _GEN_7617; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_uopc = _T_995 ? issue_slots_19_uop_uopc : _GEN_7616; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_inst = _T_995 ? issue_slots_19_uop_inst : _GEN_7615; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_inst = _T_995 ? issue_slots_19_uop_debug_inst : _GEN_7614; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_rvc = _T_995 ? issue_slots_19_uop_is_rvc : _GEN_7613; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_pc = _T_995 ? issue_slots_19_uop_debug_pc : _GEN_7612; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iq_type = _T_995 ? issue_slots_19_uop_iq_type : _GEN_7611; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_fu_code = _T_995 ? issue_slots_19_uop_fu_code : _GEN_7610; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_br_type = _T_995 ? issue_slots_19_uop_ctrl_br_type : _GEN_7609; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op1_sel = _T_995 ? issue_slots_19_uop_ctrl_op1_sel : _GEN_7608; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op2_sel = _T_995 ? issue_slots_19_uop_ctrl_op2_sel : _GEN_7607; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_imm_sel = _T_995 ? issue_slots_19_uop_ctrl_imm_sel : _GEN_7606; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op_fcn = _T_995 ? issue_slots_19_uop_ctrl_op_fcn : _GEN_7605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_fcn_dw = _T_995 ? issue_slots_19_uop_ctrl_fcn_dw : _GEN_7604; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_csr_cmd = _T_995 ? issue_slots_19_uop_ctrl_csr_cmd : _GEN_7603; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_is_load = _T_995 ? issue_slots_19_uop_ctrl_is_load : _GEN_7602; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_is_sta = _T_995 ? issue_slots_19_uop_ctrl_is_sta : _GEN_7601; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_is_std = _T_995 ? issue_slots_19_uop_ctrl_is_std : _GEN_7600; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op3_sel = _T_995 ? issue_slots_19_uop_ctrl_op3_sel : _GEN_7599; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iw_state = _T_995 ? issue_slots_19_uop_iw_state : _GEN_7598; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iw_p1_poisoned = _T_995 ? issue_slots_19_uop_iw_p1_poisoned : _GEN_7597; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iw_p2_poisoned = _T_995 ? issue_slots_19_uop_iw_p2_poisoned : _GEN_7596; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_br = _T_995 ? issue_slots_19_uop_is_br : _GEN_7595; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_jalr = _T_995 ? issue_slots_19_uop_is_jalr : _GEN_7594; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_jal = _T_995 ? issue_slots_19_uop_is_jal : _GEN_7593; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_sfb = _T_995 ? issue_slots_19_uop_is_sfb : _GEN_7592; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_br_mask = _T_995 ? issue_slots_19_uop_br_mask : _GEN_7591; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_br_tag = _T_995 ? issue_slots_19_uop_br_tag : _GEN_7590; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ftq_idx = _T_995 ? issue_slots_19_uop_ftq_idx : _GEN_7589; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_edge_inst = _T_995 ? issue_slots_19_uop_edge_inst : _GEN_7588; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pc_lob = _T_995 ? issue_slots_19_uop_pc_lob : _GEN_7587; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_taken = _T_995 ? issue_slots_19_uop_taken : _GEN_7586; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_imm_packed = _T_995 ? issue_slots_19_uop_imm_packed : _GEN_7585; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_csr_addr = _T_995 ? issue_slots_19_uop_csr_addr : _GEN_7584; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rob_idx = _T_995 ? issue_slots_19_uop_rob_idx : _GEN_7583; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldq_idx = _T_995 ? issue_slots_19_uop_ldq_idx : _GEN_7582; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_stq_idx = _T_995 ? issue_slots_19_uop_stq_idx : _GEN_7581; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rxq_idx = _T_995 ? issue_slots_19_uop_rxq_idx : _GEN_7580; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pdst = _T_995 ? issue_slots_19_uop_pdst : _GEN_7579; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs1 = _T_995 ? issue_slots_19_uop_prs1 : _GEN_7578; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs2 = _T_995 ? issue_slots_19_uop_prs2 : _GEN_7577; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs3 = _T_995 ? issue_slots_19_uop_prs3 : _GEN_7576; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ppred = _T_995 ? issue_slots_19_uop_ppred : _GEN_7575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs1_busy = _T_995 ? issue_slots_19_uop_prs1_busy : _GEN_7574; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs2_busy = _T_995 ? issue_slots_19_uop_prs2_busy : _GEN_7573; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs3_busy = _T_995 ? issue_slots_19_uop_prs3_busy : _GEN_7572; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ppred_busy = _T_995 ? issue_slots_19_uop_ppred_busy : _GEN_7571; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_stale_pdst = _T_995 ? issue_slots_19_uop_stale_pdst : _GEN_7570; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_exception = _T_995 ? issue_slots_19_uop_exception : _GEN_7569; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_exc_cause = _T_995 ? issue_slots_19_uop_exc_cause : _GEN_7568; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_bypassable = _T_995 ? issue_slots_19_uop_bypassable : _GEN_7567; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_mem_cmd = _T_995 ? issue_slots_19_uop_mem_cmd : _GEN_7566; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_mem_size = _T_995 ? issue_slots_19_uop_mem_size : _GEN_7565; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_mem_signed = _T_995 ? issue_slots_19_uop_mem_signed : _GEN_7564; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_fence = _T_995 ? issue_slots_19_uop_is_fence : _GEN_7563; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_fencei = _T_995 ? issue_slots_19_uop_is_fencei : _GEN_7562; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_amo = _T_995 ? issue_slots_19_uop_is_amo : _GEN_7561; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_uses_ldq = _T_995 ? issue_slots_19_uop_uses_ldq : _GEN_7560; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_uses_stq = _T_995 ? issue_slots_19_uop_uses_stq : _GEN_7559; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_sys_pc2epc = _T_995 ? issue_slots_19_uop_is_sys_pc2epc : _GEN_7558; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_unique = _T_995 ? issue_slots_19_uop_is_unique : _GEN_7557; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_flush_on_commit = _T_995 ? issue_slots_19_uop_flush_on_commit : _GEN_7556; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldst_is_rs1 = _T_995 ? issue_slots_19_uop_ldst_is_rs1 : _GEN_7555; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldst = _T_995 ? issue_slots_19_uop_ldst : _GEN_7554; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs1 = _T_995 ? issue_slots_19_uop_lrs1 : _GEN_7553; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs2 = _T_995 ? issue_slots_19_uop_lrs2 : _GEN_7552; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs3 = _T_995 ? issue_slots_19_uop_lrs3 : _GEN_7551; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldst_val = _T_995 ? issue_slots_19_uop_ldst_val : _GEN_7550; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_dst_rtype = _T_995 ? issue_slots_19_uop_dst_rtype : _GEN_7549; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs1_rtype = _T_995 ? issue_slots_19_uop_lrs1_rtype : _GEN_7548; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs2_rtype = _T_995 ? issue_slots_19_uop_lrs2_rtype : _GEN_7547; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_frs3_en = _T_995 ? issue_slots_19_uop_frs3_en : _GEN_7546; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_fp_val = _T_995 ? issue_slots_19_uop_fp_val : _GEN_7545; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_fp_single = _T_995 ? issue_slots_19_uop_fp_single : _GEN_7544; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_xcpt_pf_if = _T_995 ? issue_slots_19_uop_xcpt_pf_if : _GEN_7543; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_xcpt_ae_if = _T_995 ? issue_slots_19_uop_xcpt_ae_if : _GEN_7542; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_xcpt_ma_if = _T_995 ? issue_slots_19_uop_xcpt_ma_if : _GEN_7541; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_bp_debug_if = _T_995 ? issue_slots_19_uop_bp_debug_if : _GEN_7540; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_bp_xcpt_if = _T_995 ? issue_slots_19_uop_bp_xcpt_if : _GEN_7539; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_fsrc = _T_995 ? issue_slots_19_uop_debug_fsrc : _GEN_7538; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_tsrc = _T_995 ? issue_slots_19_uop_debug_tsrc : _GEN_7537; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_switch = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_switch :
    _GEN_7732; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_switch_off = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_switch_off
     : _GEN_7731; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_unicore = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_unicore
     : _GEN_7730; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_shift = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_shift :
    _GEN_7729; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_lrs3_rtype = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_lrs3_rtype
     : _GEN_7728; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_rflag = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_rflag :
    _GEN_7727; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_wflag = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_wflag :
    _GEN_7726; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_prflag = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_prflag :
    _GEN_7725; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_pwflag = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_pwflag :
    _GEN_7724; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_pflag_busy = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_pflag_busy
     : _GEN_7723; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_stale_pflag = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_stale_pflag : _GEN_7722; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_op1_sel = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_op1_sel :
    _GEN_7721; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_op2_sel = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_op2_sel :
    _GEN_7720; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_split_num = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_split_num :
    _GEN_7719; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_self_index = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_self_index
     : _GEN_7718; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_rob_inst_idx = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_rob_inst_idx : _GEN_7717; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_address_num = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_address_num : _GEN_7716; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_uopc = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_uopc : _GEN_7715; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_inst = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_inst : _GEN_7714; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_debug_inst = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_debug_inst
     : _GEN_7713; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_rvc = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_rvc :
    _GEN_7712; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_debug_pc = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_debug_pc :
    _GEN_7711; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_iq_type = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_iq_type :
    _GEN_7710; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_fu_code = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_fu_code :
    _GEN_7709; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_br_type = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_br_type : _GEN_7708; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_op1_sel = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_op1_sel : _GEN_7707; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_op2_sel = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_op2_sel : _GEN_7706; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_imm_sel = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_imm_sel : _GEN_7705; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_op_fcn = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_op_fcn : _GEN_7704; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_fcn_dw = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_fcn_dw : _GEN_7703; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_csr_cmd = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_csr_cmd : _GEN_7702; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_is_load = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_is_load : _GEN_7701; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_is_sta = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_is_sta : _GEN_7700; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_is_std = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_is_std : _GEN_7699; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ctrl_op3_sel = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ctrl_op3_sel : _GEN_7698; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_iw_state = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_iw_state :
    _GEN_7697; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_iw_p1_poisoned = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_iw_p1_poisoned : _GEN_7696; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_iw_p2_poisoned = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_iw_p2_poisoned : _GEN_7695; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_br = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_br :
    _GEN_7694; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_jalr = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_jalr :
    _GEN_7693; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_jal = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_jal :
    _GEN_7692; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_sfb = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_sfb :
    _GEN_7691; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_br_mask = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_br_mask :
    _GEN_7690; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_br_tag = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_br_tag :
    _GEN_7689; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ftq_idx = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_ftq_idx :
    _GEN_7688; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_edge_inst = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_edge_inst :
    _GEN_7687; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_pc_lob = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_pc_lob :
    _GEN_7686; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_taken = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_taken :
    _GEN_7685; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_imm_packed = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_imm_packed
     : _GEN_7684; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_csr_addr = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_csr_addr :
    _GEN_7683; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_rob_idx = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_rob_idx :
    _GEN_7682; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ldq_idx = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_ldq_idx :
    _GEN_7681; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_stq_idx = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_stq_idx :
    _GEN_7680; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_rxq_idx = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_rxq_idx :
    _GEN_7679; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_pdst = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_pdst : _GEN_7678; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_prs1 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_prs1 : _GEN_7677; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_prs2 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_prs2 : _GEN_7676; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_prs3 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_prs3 : _GEN_7675; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ppred = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_ppred :
    _GEN_7674; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_prs1_busy = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_prs1_busy :
    _GEN_7673; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_prs2_busy = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_prs2_busy :
    _GEN_7672; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_prs3_busy = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_prs3_busy :
    _GEN_7671; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ppred_busy = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_ppred_busy
     : _GEN_7670; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_stale_pdst = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_stale_pdst
     : _GEN_7669; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_exception = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_exception :
    _GEN_7668; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_exc_cause = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_exc_cause :
    _GEN_7667; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_bypassable = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_bypassable
     : _GEN_7666; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_mem_cmd = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_mem_cmd :
    _GEN_7665; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_mem_size = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_mem_size :
    _GEN_7664; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_mem_signed = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_mem_signed
     : _GEN_7663; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_fence = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_fence :
    _GEN_7662; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_fencei = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_fencei :
    _GEN_7661; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_amo = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_amo :
    _GEN_7660; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_uses_ldq = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_uses_ldq :
    _GEN_7659; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_uses_stq = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_uses_stq :
    _GEN_7658; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_sys_pc2epc = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_is_sys_pc2epc : _GEN_7657; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_is_unique = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_is_unique :
    _GEN_7656; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_flush_on_commit = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_flush_on_commit : _GEN_7655; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ldst_is_rs1 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_ldst_is_rs1 : _GEN_7654; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ldst = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_ldst : _GEN_7653; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_lrs1 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_lrs1 : _GEN_7652; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_lrs2 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_lrs2 : _GEN_7651; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_lrs3 = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_lrs3 : _GEN_7650; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_ldst_val = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_ldst_val :
    _GEN_7649; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_dst_rtype = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_dst_rtype :
    _GEN_7648; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_lrs1_rtype = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_lrs1_rtype
     : _GEN_7647; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_lrs2_rtype = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_lrs2_rtype
     : _GEN_7646; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_frs3_en = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_frs3_en :
    _GEN_7645; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_fp_val = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_fp_val :
    _GEN_7644; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_fp_single = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_fp_single :
    _GEN_7643; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_xcpt_pf_if = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_xcpt_pf_if
     : _GEN_7642; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_xcpt_ae_if = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_xcpt_ae_if
     : _GEN_7641; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_xcpt_ma_if = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_xcpt_ma_if
     : _GEN_7640; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_bp_debug_if = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ?
    issue_slots_19_uop_bp_debug_if : _GEN_7639; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_bp_xcpt_if = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_bp_xcpt_if
     : _GEN_7638; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_debug_fsrc = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_debug_fsrc
     : _GEN_7637; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_1_debug_tsrc = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 ? issue_slots_19_uop_debug_tsrc
     : _GEN_7636; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_event_empty = ~(issue_slots_0_valid | issue_slots_1_valid | issue_slots_2_valid | issue_slots_3_valid |
    issue_slots_4_valid | issue_slots_5_valid | issue_slots_6_valid | issue_slots_7_valid | issue_slots_8_valid |
    issue_slots_9_valid | issue_slots_10_valid | issue_slots_11_valid | issue_slots_12_valid | issue_slots_13_valid |
    issue_slots_14_valid | issue_slots_15_valid | issue_slots_16_valid | issue_slots_17_valid | issue_slots_18_valid |
    issue_slots_19_valid); // @[issue-unit.scala 169:21]
  assign slots_0_clock = clock;
  assign slots_0_reset = reset;
  assign slots_0_io_grant = issue_slots_0_request & ~_T_423 & _T_428 | _T_423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_0_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_0_io_clear = 1'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_0_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_0_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_0_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_0_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_0_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_0_io_in_uop_valid = _GEN_13[1:0] == 2'h2 ? issue_slots_2_will_be_valid : _GEN_52; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_0_io_in_uop_bits_switch = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_switch :
    issue_slots_1_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_switch_off = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_switch_off :
    issue_slots_1_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_unicore = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_unicore :
    issue_slots_1_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_shift = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_shift : issue_slots_1_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs3_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs3_rtype :
    issue_slots_1_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rflag = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_rflag : issue_slots_1_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_wflag = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_wflag : issue_slots_1_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prflag = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prflag :
    issue_slots_1_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pwflag = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_pwflag :
    issue_slots_1_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pflag_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_pflag_busy :
    issue_slots_1_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stale_pflag = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_stale_pflag :
    issue_slots_1_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_op1_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_op1_sel :
    issue_slots_1_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_op2_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_op2_sel :
    issue_slots_1_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_split_num = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_split_num :
    issue_slots_1_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_self_index = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_self_index :
    issue_slots_1_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rob_inst_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_rob_inst_idx :
    issue_slots_1_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_address_num = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_address_num :
    issue_slots_1_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uopc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_uopc : issue_slots_1_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_inst : issue_slots_1_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_inst :
    issue_slots_1_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_rvc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_rvc :
    issue_slots_1_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_pc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_pc :
    issue_slots_1_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iq_type = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iq_type :
    issue_slots_1_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fu_code = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_fu_code :
    issue_slots_1_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_br_type = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_br_type :
    issue_slots_1_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op1_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op1_sel :
    issue_slots_1_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op2_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op2_sel :
    issue_slots_1_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_imm_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_imm_sel :
    issue_slots_1_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op_fcn = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op_fcn :
    issue_slots_1_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_fcn_dw = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_fcn_dw :
    issue_slots_1_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_csr_cmd = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_csr_cmd :
    issue_slots_1_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_load = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_load :
    issue_slots_1_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_sta = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_sta :
    issue_slots_1_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_std = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_std :
    issue_slots_1_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op3_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op3_sel :
    issue_slots_1_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_state = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_state :
    issue_slots_1_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_p1_poisoned = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_p1_poisoned :
    issue_slots_1_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_p2_poisoned = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_p2_poisoned :
    issue_slots_1_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_br = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_br : issue_slots_1_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_jalr = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_jalr :
    issue_slots_1_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_jal = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_jal :
    issue_slots_1_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_sfb = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_sfb :
    issue_slots_1_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_br_mask = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_br_mask :
    issue_slots_1_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_br_tag = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_br_tag :
    issue_slots_1_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ftq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ftq_idx :
    issue_slots_1_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_edge_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_edge_inst :
    issue_slots_1_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pc_lob = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_pc_lob :
    issue_slots_1_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_taken = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_taken : issue_slots_1_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_imm_packed = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_imm_packed :
    issue_slots_1_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_csr_addr = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_csr_addr :
    issue_slots_1_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rob_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_rob_idx :
    issue_slots_1_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldq_idx :
    issue_slots_1_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_stq_idx :
    issue_slots_1_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rxq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_rxq_idx :
    issue_slots_1_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pdst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_pdst : issue_slots_1_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs1 : issue_slots_1_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs2 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs2 : issue_slots_1_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs3 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs3 : issue_slots_1_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ppred = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ppred : issue_slots_1_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs1_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs1_busy :
    issue_slots_1_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs2_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs2_busy :
    issue_slots_1_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs3_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs3_busy :
    issue_slots_1_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ppred_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ppred_busy :
    issue_slots_1_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stale_pdst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_stale_pdst :
    issue_slots_1_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_exception = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_exception :
    issue_slots_1_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_exc_cause = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_exc_cause :
    issue_slots_1_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bypassable = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_bypassable :
    issue_slots_1_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_cmd = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_cmd :
    issue_slots_1_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_size = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_size :
    issue_slots_1_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_signed = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_signed :
    issue_slots_1_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_fence = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_fence :
    issue_slots_1_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_fencei = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_fencei :
    issue_slots_1_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_amo = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_amo :
    issue_slots_1_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uses_ldq = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_uses_ldq :
    issue_slots_1_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uses_stq = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_uses_stq :
    issue_slots_1_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_sys_pc2epc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_sys_pc2epc :
    issue_slots_1_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_unique = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_unique :
    issue_slots_1_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_flush_on_commit = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_flush_on_commit :
    issue_slots_1_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst_is_rs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst_is_rs1 :
    issue_slots_1_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst : issue_slots_1_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs1 : issue_slots_1_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs2 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs2 : issue_slots_1_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs3 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs3 : issue_slots_1_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst_val = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst_val :
    issue_slots_1_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_dst_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_dst_rtype :
    issue_slots_1_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs1_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs1_rtype :
    issue_slots_1_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs2_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs2_rtype :
    issue_slots_1_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_frs3_en = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_frs3_en :
    issue_slots_1_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fp_val = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_fp_val :
    issue_slots_1_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fp_single = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_fp_single :
    issue_slots_1_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_pf_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_pf_if :
    issue_slots_1_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_ae_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_ae_if :
    issue_slots_1_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_ma_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_ma_if :
    issue_slots_1_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bp_debug_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_bp_debug_if :
    issue_slots_1_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bp_xcpt_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_bp_xcpt_if :
    issue_slots_1_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_fsrc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_fsrc :
    issue_slots_1_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_tsrc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_tsrc :
    issue_slots_1_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_clock = clock;
  assign slots_1_reset = reset;
  assign slots_1_io_grant = issue_slots_1_request & ~_T_455 & _T_458 & ~(issue_slots_0_request & ~_T_423 & _T_428) |
    _T_455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_1_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_1_io_clear = _GEN_11[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_1_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_1_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_1_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_1_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_1_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_1_io_in_uop_valid = _GEN_15[1:0] == 2'h2 ? issue_slots_3_will_be_valid : _GEN_248; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_1_io_in_uop_bits_switch = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_switch :
    issue_slots_2_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_switch_off = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_switch_off :
    issue_slots_2_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_unicore = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_unicore :
    issue_slots_2_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_shift = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_shift : issue_slots_2_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs3_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs3_rtype :
    issue_slots_2_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rflag = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_rflag : issue_slots_2_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_wflag = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_wflag : issue_slots_2_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prflag = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prflag :
    issue_slots_2_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pwflag = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_pwflag :
    issue_slots_2_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pflag_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_pflag_busy :
    issue_slots_2_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stale_pflag = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_stale_pflag :
    issue_slots_2_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_op1_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_op1_sel :
    issue_slots_2_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_op2_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_op2_sel :
    issue_slots_2_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_split_num = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_split_num :
    issue_slots_2_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_self_index = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_self_index :
    issue_slots_2_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rob_inst_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_rob_inst_idx :
    issue_slots_2_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_address_num = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_address_num :
    issue_slots_2_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uopc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_uopc : issue_slots_2_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_inst : issue_slots_2_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_inst :
    issue_slots_2_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_rvc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_rvc :
    issue_slots_2_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_pc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_pc :
    issue_slots_2_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iq_type = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iq_type :
    issue_slots_2_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fu_code = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_fu_code :
    issue_slots_2_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_br_type = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_br_type :
    issue_slots_2_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op1_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op1_sel :
    issue_slots_2_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op2_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op2_sel :
    issue_slots_2_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_imm_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_imm_sel :
    issue_slots_2_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op_fcn = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op_fcn :
    issue_slots_2_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_fcn_dw = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_fcn_dw :
    issue_slots_2_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_csr_cmd = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_csr_cmd :
    issue_slots_2_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_load = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_load :
    issue_slots_2_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_sta = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_sta :
    issue_slots_2_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_std = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_std :
    issue_slots_2_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op3_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op3_sel :
    issue_slots_2_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_state = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_state :
    issue_slots_2_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_p1_poisoned = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_p1_poisoned :
    issue_slots_2_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_p2_poisoned = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_p2_poisoned :
    issue_slots_2_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_br = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_br : issue_slots_2_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_jalr = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_jalr :
    issue_slots_2_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_jal = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_jal :
    issue_slots_2_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_sfb = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_sfb :
    issue_slots_2_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_br_mask = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_br_mask :
    issue_slots_2_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_br_tag = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_br_tag :
    issue_slots_2_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ftq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ftq_idx :
    issue_slots_2_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_edge_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_edge_inst :
    issue_slots_2_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pc_lob = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_pc_lob :
    issue_slots_2_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_taken = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_taken : issue_slots_2_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_imm_packed = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_imm_packed :
    issue_slots_2_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_csr_addr = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_csr_addr :
    issue_slots_2_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rob_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_rob_idx :
    issue_slots_2_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldq_idx :
    issue_slots_2_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_stq_idx :
    issue_slots_2_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rxq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_rxq_idx :
    issue_slots_2_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pdst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_pdst : issue_slots_2_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs1 : issue_slots_2_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs2 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs2 : issue_slots_2_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs3 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs3 : issue_slots_2_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ppred = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ppred : issue_slots_2_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs1_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs1_busy :
    issue_slots_2_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs2_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs2_busy :
    issue_slots_2_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs3_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs3_busy :
    issue_slots_2_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ppred_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ppred_busy :
    issue_slots_2_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stale_pdst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_stale_pdst :
    issue_slots_2_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_exception = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_exception :
    issue_slots_2_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_exc_cause = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_exc_cause :
    issue_slots_2_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bypassable = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_bypassable :
    issue_slots_2_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_cmd = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_cmd :
    issue_slots_2_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_size = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_size :
    issue_slots_2_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_signed = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_signed :
    issue_slots_2_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_fence = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_fence :
    issue_slots_2_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_fencei = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_fencei :
    issue_slots_2_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_amo = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_amo :
    issue_slots_2_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uses_ldq = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_uses_ldq :
    issue_slots_2_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uses_stq = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_uses_stq :
    issue_slots_2_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_sys_pc2epc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_sys_pc2epc :
    issue_slots_2_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_unique = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_unique :
    issue_slots_2_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_flush_on_commit = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_flush_on_commit :
    issue_slots_2_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst_is_rs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst_is_rs1 :
    issue_slots_2_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst : issue_slots_2_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs1 : issue_slots_2_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs2 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs2 : issue_slots_2_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs3 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs3 : issue_slots_2_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst_val = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst_val :
    issue_slots_2_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_dst_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_dst_rtype :
    issue_slots_2_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs1_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs1_rtype :
    issue_slots_2_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs2_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs2_rtype :
    issue_slots_2_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_frs3_en = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_frs3_en :
    issue_slots_2_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fp_val = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_fp_val :
    issue_slots_2_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fp_single = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_fp_single :
    issue_slots_2_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_pf_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_pf_if :
    issue_slots_2_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_ae_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_ae_if :
    issue_slots_2_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_ma_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_ma_if :
    issue_slots_2_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bp_debug_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_bp_debug_if :
    issue_slots_2_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bp_xcpt_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_bp_xcpt_if :
    issue_slots_2_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_fsrc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_fsrc :
    issue_slots_2_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_tsrc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_tsrc :
    issue_slots_2_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_clock = clock;
  assign slots_2_reset = reset;
  assign slots_2_io_grant = _T_496 & ~_T_467 | _T_485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_2_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_2_io_clear = _GEN_13[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_2_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_2_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_2_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_2_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_2_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_2_io_in_uop_valid = _GEN_17[1:0] == 2'h2 ? issue_slots_4_will_be_valid : _GEN_444; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_2_io_in_uop_bits_switch = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_switch :
    issue_slots_3_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_switch_off = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_switch_off :
    issue_slots_3_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_unicore = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_unicore :
    issue_slots_3_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_shift = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_shift : issue_slots_3_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs3_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs3_rtype :
    issue_slots_3_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rflag = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_rflag : issue_slots_3_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_wflag = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_wflag : issue_slots_3_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prflag = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prflag :
    issue_slots_3_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pwflag = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_pwflag :
    issue_slots_3_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pflag_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_pflag_busy :
    issue_slots_3_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stale_pflag = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_stale_pflag :
    issue_slots_3_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_op1_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_op1_sel :
    issue_slots_3_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_op2_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_op2_sel :
    issue_slots_3_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_split_num = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_split_num :
    issue_slots_3_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_self_index = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_self_index :
    issue_slots_3_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rob_inst_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_rob_inst_idx :
    issue_slots_3_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_address_num = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_address_num :
    issue_slots_3_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uopc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_uopc : issue_slots_3_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_inst : issue_slots_3_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_inst :
    issue_slots_3_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_rvc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_rvc :
    issue_slots_3_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_pc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_pc :
    issue_slots_3_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iq_type = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iq_type :
    issue_slots_3_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fu_code = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_fu_code :
    issue_slots_3_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_br_type = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_br_type :
    issue_slots_3_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op1_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op1_sel :
    issue_slots_3_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op2_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op2_sel :
    issue_slots_3_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_imm_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_imm_sel :
    issue_slots_3_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op_fcn = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op_fcn :
    issue_slots_3_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_fcn_dw = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_fcn_dw :
    issue_slots_3_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_csr_cmd = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_csr_cmd :
    issue_slots_3_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_load = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_load :
    issue_slots_3_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_sta = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_sta :
    issue_slots_3_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_std = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_std :
    issue_slots_3_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op3_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op3_sel :
    issue_slots_3_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_state = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_state :
    issue_slots_3_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_p1_poisoned = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_p1_poisoned :
    issue_slots_3_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_p2_poisoned = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_p2_poisoned :
    issue_slots_3_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_br = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_br : issue_slots_3_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_jalr = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_jalr :
    issue_slots_3_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_jal = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_jal :
    issue_slots_3_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_sfb = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_sfb :
    issue_slots_3_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_br_mask = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_br_mask :
    issue_slots_3_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_br_tag = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_br_tag :
    issue_slots_3_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ftq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ftq_idx :
    issue_slots_3_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_edge_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_edge_inst :
    issue_slots_3_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pc_lob = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_pc_lob :
    issue_slots_3_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_taken = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_taken : issue_slots_3_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_imm_packed = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_imm_packed :
    issue_slots_3_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_csr_addr = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_csr_addr :
    issue_slots_3_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rob_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_rob_idx :
    issue_slots_3_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldq_idx :
    issue_slots_3_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_stq_idx :
    issue_slots_3_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rxq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_rxq_idx :
    issue_slots_3_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pdst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_pdst : issue_slots_3_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs1 : issue_slots_3_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs2 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs2 : issue_slots_3_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs3 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs3 : issue_slots_3_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ppred = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ppred : issue_slots_3_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs1_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs1_busy :
    issue_slots_3_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs2_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs2_busy :
    issue_slots_3_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs3_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs3_busy :
    issue_slots_3_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ppred_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ppred_busy :
    issue_slots_3_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stale_pdst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_stale_pdst :
    issue_slots_3_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_exception = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_exception :
    issue_slots_3_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_exc_cause = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_exc_cause :
    issue_slots_3_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bypassable = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_bypassable :
    issue_slots_3_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_cmd = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_cmd :
    issue_slots_3_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_size = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_size :
    issue_slots_3_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_signed = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_signed :
    issue_slots_3_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_fence = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_fence :
    issue_slots_3_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_fencei = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_fencei :
    issue_slots_3_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_amo = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_amo :
    issue_slots_3_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uses_ldq = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_uses_ldq :
    issue_slots_3_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uses_stq = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_uses_stq :
    issue_slots_3_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_sys_pc2epc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_sys_pc2epc :
    issue_slots_3_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_unique = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_unique :
    issue_slots_3_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_flush_on_commit = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_flush_on_commit :
    issue_slots_3_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst_is_rs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst_is_rs1 :
    issue_slots_3_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst : issue_slots_3_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs1 : issue_slots_3_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs2 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs2 : issue_slots_3_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs3 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs3 : issue_slots_3_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst_val = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst_val :
    issue_slots_3_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_dst_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_dst_rtype :
    issue_slots_3_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs1_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs1_rtype :
    issue_slots_3_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs2_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs2_rtype :
    issue_slots_3_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_frs3_en = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_frs3_en :
    issue_slots_3_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fp_val = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_fp_val :
    issue_slots_3_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fp_single = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_fp_single :
    issue_slots_3_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_pf_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_pf_if :
    issue_slots_3_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_ae_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_ae_if :
    issue_slots_3_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_ma_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_ma_if :
    issue_slots_3_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bp_debug_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_bp_debug_if :
    issue_slots_3_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bp_xcpt_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_bp_xcpt_if :
    issue_slots_3_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_fsrc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_fsrc :
    issue_slots_3_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_tsrc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_tsrc :
    issue_slots_3_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_clock = clock;
  assign slots_3_reset = reset;
  assign slots_3_io_grant = issue_slots_3_request & ~_T_515 & _T_518 & ~_T_497 | _T_515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_3_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_3_io_clear = _GEN_15[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_3_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_3_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_3_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_3_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_3_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_3_io_in_uop_valid = _GEN_19[1:0] == 2'h2 ? issue_slots_5_will_be_valid : _GEN_640; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_3_io_in_uop_bits_switch = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_switch :
    issue_slots_4_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_switch_off = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_switch_off :
    issue_slots_4_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_unicore = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_unicore :
    issue_slots_4_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_shift = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_shift : issue_slots_4_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs3_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs3_rtype :
    issue_slots_4_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rflag = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_rflag : issue_slots_4_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_wflag = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_wflag : issue_slots_4_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prflag = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prflag :
    issue_slots_4_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pwflag = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_pwflag :
    issue_slots_4_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pflag_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_pflag_busy :
    issue_slots_4_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stale_pflag = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_stale_pflag :
    issue_slots_4_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_op1_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_op1_sel :
    issue_slots_4_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_op2_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_op2_sel :
    issue_slots_4_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_split_num = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_split_num :
    issue_slots_4_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_self_index = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_self_index :
    issue_slots_4_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rob_inst_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_rob_inst_idx :
    issue_slots_4_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_address_num = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_address_num :
    issue_slots_4_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uopc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_uopc : issue_slots_4_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_inst : issue_slots_4_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_inst :
    issue_slots_4_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_rvc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_rvc :
    issue_slots_4_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_pc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_pc :
    issue_slots_4_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iq_type = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iq_type :
    issue_slots_4_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fu_code = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_fu_code :
    issue_slots_4_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_br_type = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_br_type :
    issue_slots_4_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op1_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op1_sel :
    issue_slots_4_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op2_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op2_sel :
    issue_slots_4_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_imm_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_imm_sel :
    issue_slots_4_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op_fcn = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op_fcn :
    issue_slots_4_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_fcn_dw = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_fcn_dw :
    issue_slots_4_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_csr_cmd = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_csr_cmd :
    issue_slots_4_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_load = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_load :
    issue_slots_4_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_sta = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_sta :
    issue_slots_4_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_std = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_std :
    issue_slots_4_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op3_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op3_sel :
    issue_slots_4_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_state = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_state :
    issue_slots_4_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_p1_poisoned = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_p1_poisoned :
    issue_slots_4_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_p2_poisoned = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_p2_poisoned :
    issue_slots_4_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_br = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_br : issue_slots_4_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_jalr = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_jalr :
    issue_slots_4_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_jal = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_jal :
    issue_slots_4_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_sfb = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_sfb :
    issue_slots_4_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_br_mask = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_br_mask :
    issue_slots_4_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_br_tag = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_br_tag :
    issue_slots_4_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ftq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ftq_idx :
    issue_slots_4_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_edge_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_edge_inst :
    issue_slots_4_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pc_lob = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_pc_lob :
    issue_slots_4_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_taken = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_taken : issue_slots_4_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_imm_packed = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_imm_packed :
    issue_slots_4_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_csr_addr = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_csr_addr :
    issue_slots_4_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rob_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_rob_idx :
    issue_slots_4_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldq_idx :
    issue_slots_4_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_stq_idx :
    issue_slots_4_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rxq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_rxq_idx :
    issue_slots_4_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pdst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_pdst : issue_slots_4_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs1 : issue_slots_4_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs2 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs2 : issue_slots_4_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs3 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs3 : issue_slots_4_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ppred = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ppred : issue_slots_4_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs1_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs1_busy :
    issue_slots_4_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs2_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs2_busy :
    issue_slots_4_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs3_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs3_busy :
    issue_slots_4_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ppred_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ppred_busy :
    issue_slots_4_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stale_pdst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_stale_pdst :
    issue_slots_4_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_exception = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_exception :
    issue_slots_4_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_exc_cause = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_exc_cause :
    issue_slots_4_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bypassable = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_bypassable :
    issue_slots_4_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_cmd = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_cmd :
    issue_slots_4_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_size = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_size :
    issue_slots_4_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_signed = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_signed :
    issue_slots_4_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_fence = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_fence :
    issue_slots_4_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_fencei = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_fencei :
    issue_slots_4_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_amo = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_amo :
    issue_slots_4_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uses_ldq = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_uses_ldq :
    issue_slots_4_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uses_stq = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_uses_stq :
    issue_slots_4_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_sys_pc2epc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_sys_pc2epc :
    issue_slots_4_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_unique = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_unique :
    issue_slots_4_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_flush_on_commit = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_flush_on_commit :
    issue_slots_4_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst_is_rs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst_is_rs1 :
    issue_slots_4_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst : issue_slots_4_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs1 : issue_slots_4_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs2 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs2 : issue_slots_4_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs3 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs3 : issue_slots_4_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst_val = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst_val :
    issue_slots_4_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_dst_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_dst_rtype :
    issue_slots_4_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs1_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs1_rtype :
    issue_slots_4_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs2_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs2_rtype :
    issue_slots_4_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_frs3_en = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_frs3_en :
    issue_slots_4_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fp_val = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_fp_val :
    issue_slots_4_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fp_single = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_fp_single :
    issue_slots_4_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_pf_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_pf_if :
    issue_slots_4_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_ae_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_ae_if :
    issue_slots_4_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_ma_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_ma_if :
    issue_slots_4_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bp_debug_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_bp_debug_if :
    issue_slots_4_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bp_xcpt_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_bp_xcpt_if :
    issue_slots_4_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_fsrc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_fsrc :
    issue_slots_4_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_tsrc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_tsrc :
    issue_slots_4_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_clock = clock;
  assign slots_4_reset = reset;
  assign slots_4_io_grant = issue_slots_4_request & ~_T_545 & _T_548 & ~_T_527 | _T_545; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_4_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_4_io_clear = _GEN_17[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_4_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_4_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_4_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_4_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_4_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_4_io_in_uop_valid = _GEN_21[1:0] == 2'h2 ? issue_slots_6_will_be_valid : _GEN_836; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_4_io_in_uop_bits_switch = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_switch :
    issue_slots_5_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_switch_off = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_switch_off :
    issue_slots_5_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_unicore = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_unicore :
    issue_slots_5_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_shift = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_shift : issue_slots_5_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs3_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs3_rtype :
    issue_slots_5_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rflag = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_rflag : issue_slots_5_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_wflag = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_wflag : issue_slots_5_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prflag = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prflag :
    issue_slots_5_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pwflag = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_pwflag :
    issue_slots_5_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pflag_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_pflag_busy :
    issue_slots_5_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stale_pflag = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_stale_pflag :
    issue_slots_5_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_op1_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_op1_sel :
    issue_slots_5_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_op2_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_op2_sel :
    issue_slots_5_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_split_num = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_split_num :
    issue_slots_5_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_self_index = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_self_index :
    issue_slots_5_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rob_inst_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_rob_inst_idx :
    issue_slots_5_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_address_num = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_address_num :
    issue_slots_5_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uopc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_uopc : issue_slots_5_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_inst : issue_slots_5_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_inst :
    issue_slots_5_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_rvc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_rvc :
    issue_slots_5_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_pc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_pc :
    issue_slots_5_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iq_type = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iq_type :
    issue_slots_5_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fu_code = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_fu_code :
    issue_slots_5_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_br_type = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_br_type :
    issue_slots_5_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op1_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op1_sel :
    issue_slots_5_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op2_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op2_sel :
    issue_slots_5_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_imm_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_imm_sel :
    issue_slots_5_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op_fcn = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op_fcn :
    issue_slots_5_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_fcn_dw = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_fcn_dw :
    issue_slots_5_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_csr_cmd = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_csr_cmd :
    issue_slots_5_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_load = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_load :
    issue_slots_5_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_sta = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_sta :
    issue_slots_5_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_std = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_std :
    issue_slots_5_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op3_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op3_sel :
    issue_slots_5_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_state = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_state :
    issue_slots_5_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_p1_poisoned = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_p1_poisoned :
    issue_slots_5_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_p2_poisoned = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_p2_poisoned :
    issue_slots_5_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_br = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_br : issue_slots_5_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_jalr = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_jalr :
    issue_slots_5_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_jal = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_jal :
    issue_slots_5_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_sfb = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_sfb :
    issue_slots_5_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_br_mask = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_br_mask :
    issue_slots_5_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_br_tag = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_br_tag :
    issue_slots_5_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ftq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ftq_idx :
    issue_slots_5_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_edge_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_edge_inst :
    issue_slots_5_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pc_lob = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_pc_lob :
    issue_slots_5_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_taken = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_taken : issue_slots_5_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_imm_packed = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_imm_packed :
    issue_slots_5_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_csr_addr = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_csr_addr :
    issue_slots_5_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rob_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_rob_idx :
    issue_slots_5_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldq_idx :
    issue_slots_5_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_stq_idx :
    issue_slots_5_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rxq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_rxq_idx :
    issue_slots_5_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pdst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_pdst : issue_slots_5_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs1 : issue_slots_5_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs2 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs2 : issue_slots_5_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs3 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs3 : issue_slots_5_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ppred = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ppred : issue_slots_5_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs1_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs1_busy :
    issue_slots_5_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs2_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs2_busy :
    issue_slots_5_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs3_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs3_busy :
    issue_slots_5_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ppred_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ppred_busy :
    issue_slots_5_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stale_pdst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_stale_pdst :
    issue_slots_5_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_exception = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_exception :
    issue_slots_5_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_exc_cause = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_exc_cause :
    issue_slots_5_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bypassable = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_bypassable :
    issue_slots_5_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_cmd = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_cmd :
    issue_slots_5_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_size = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_size :
    issue_slots_5_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_signed = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_signed :
    issue_slots_5_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_fence = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_fence :
    issue_slots_5_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_fencei = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_fencei :
    issue_slots_5_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_amo = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_amo :
    issue_slots_5_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uses_ldq = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_uses_ldq :
    issue_slots_5_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uses_stq = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_uses_stq :
    issue_slots_5_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_sys_pc2epc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_sys_pc2epc :
    issue_slots_5_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_unique = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_unique :
    issue_slots_5_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_flush_on_commit = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_flush_on_commit :
    issue_slots_5_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst_is_rs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst_is_rs1 :
    issue_slots_5_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst : issue_slots_5_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs1 : issue_slots_5_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs2 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs2 : issue_slots_5_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs3 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs3 : issue_slots_5_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst_val = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst_val :
    issue_slots_5_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_dst_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_dst_rtype :
    issue_slots_5_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs1_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs1_rtype :
    issue_slots_5_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs2_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs2_rtype :
    issue_slots_5_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_frs3_en = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_frs3_en :
    issue_slots_5_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fp_val = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_fp_val :
    issue_slots_5_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fp_single = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_fp_single :
    issue_slots_5_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_pf_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_pf_if :
    issue_slots_5_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_ae_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_ae_if :
    issue_slots_5_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_ma_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_ma_if :
    issue_slots_5_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bp_debug_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_bp_debug_if :
    issue_slots_5_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bp_xcpt_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_bp_xcpt_if :
    issue_slots_5_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_fsrc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_fsrc :
    issue_slots_5_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_tsrc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_tsrc :
    issue_slots_5_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_clock = clock;
  assign slots_5_reset = reset;
  assign slots_5_io_grant = issue_slots_5_request & ~_T_575 & _T_578 & ~_T_557 | _T_575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_5_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_5_io_clear = _GEN_19[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_5_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_5_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_5_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_5_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_5_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_5_io_in_uop_valid = _GEN_23[1:0] == 2'h2 ? issue_slots_7_will_be_valid : _GEN_1032; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_5_io_in_uop_bits_switch = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_switch :
    issue_slots_6_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_switch_off = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_switch_off :
    issue_slots_6_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_unicore = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_unicore :
    issue_slots_6_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_shift = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_shift : issue_slots_6_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs3_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs3_rtype :
    issue_slots_6_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rflag = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_rflag : issue_slots_6_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_wflag = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_wflag : issue_slots_6_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prflag = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prflag :
    issue_slots_6_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pwflag = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_pwflag :
    issue_slots_6_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pflag_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_pflag_busy :
    issue_slots_6_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stale_pflag = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_stale_pflag :
    issue_slots_6_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_op1_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_op1_sel :
    issue_slots_6_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_op2_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_op2_sel :
    issue_slots_6_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_split_num = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_split_num :
    issue_slots_6_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_self_index = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_self_index :
    issue_slots_6_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rob_inst_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_rob_inst_idx :
    issue_slots_6_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_address_num = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_address_num :
    issue_slots_6_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uopc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_uopc : issue_slots_6_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_inst : issue_slots_6_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_inst :
    issue_slots_6_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_rvc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_rvc :
    issue_slots_6_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_pc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_pc :
    issue_slots_6_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iq_type = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iq_type :
    issue_slots_6_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fu_code = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_fu_code :
    issue_slots_6_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_br_type = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_br_type :
    issue_slots_6_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op1_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op1_sel :
    issue_slots_6_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op2_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op2_sel :
    issue_slots_6_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_imm_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_imm_sel :
    issue_slots_6_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op_fcn = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op_fcn :
    issue_slots_6_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_fcn_dw = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_fcn_dw :
    issue_slots_6_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_csr_cmd = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_csr_cmd :
    issue_slots_6_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_load = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_load :
    issue_slots_6_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_sta = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_sta :
    issue_slots_6_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_std = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_std :
    issue_slots_6_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op3_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op3_sel :
    issue_slots_6_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_state = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_state :
    issue_slots_6_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_p1_poisoned = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_p1_poisoned :
    issue_slots_6_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_p2_poisoned = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_p2_poisoned :
    issue_slots_6_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_br = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_br : issue_slots_6_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_jalr = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_jalr :
    issue_slots_6_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_jal = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_jal :
    issue_slots_6_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_sfb = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_sfb :
    issue_slots_6_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_br_mask = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_br_mask :
    issue_slots_6_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_br_tag = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_br_tag :
    issue_slots_6_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ftq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ftq_idx :
    issue_slots_6_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_edge_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_edge_inst :
    issue_slots_6_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pc_lob = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_pc_lob :
    issue_slots_6_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_taken = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_taken : issue_slots_6_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_imm_packed = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_imm_packed :
    issue_slots_6_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_csr_addr = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_csr_addr :
    issue_slots_6_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rob_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_rob_idx :
    issue_slots_6_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldq_idx :
    issue_slots_6_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_stq_idx :
    issue_slots_6_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rxq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_rxq_idx :
    issue_slots_6_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pdst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_pdst : issue_slots_6_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs1 : issue_slots_6_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs2 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs2 : issue_slots_6_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs3 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs3 : issue_slots_6_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ppred = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ppred : issue_slots_6_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs1_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs1_busy :
    issue_slots_6_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs2_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs2_busy :
    issue_slots_6_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs3_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs3_busy :
    issue_slots_6_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ppred_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ppred_busy :
    issue_slots_6_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stale_pdst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_stale_pdst :
    issue_slots_6_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_exception = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_exception :
    issue_slots_6_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_exc_cause = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_exc_cause :
    issue_slots_6_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bypassable = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_bypassable :
    issue_slots_6_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_cmd = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_cmd :
    issue_slots_6_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_size = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_size :
    issue_slots_6_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_signed = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_signed :
    issue_slots_6_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_fence = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_fence :
    issue_slots_6_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_fencei = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_fencei :
    issue_slots_6_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_amo = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_amo :
    issue_slots_6_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uses_ldq = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_uses_ldq :
    issue_slots_6_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uses_stq = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_uses_stq :
    issue_slots_6_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_sys_pc2epc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_sys_pc2epc :
    issue_slots_6_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_unique = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_unique :
    issue_slots_6_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_flush_on_commit = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_flush_on_commit :
    issue_slots_6_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst_is_rs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst_is_rs1 :
    issue_slots_6_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst : issue_slots_6_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs1 : issue_slots_6_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs2 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs2 : issue_slots_6_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs3 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs3 : issue_slots_6_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst_val = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst_val :
    issue_slots_6_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_dst_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_dst_rtype :
    issue_slots_6_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs1_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs1_rtype :
    issue_slots_6_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs2_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs2_rtype :
    issue_slots_6_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_frs3_en = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_frs3_en :
    issue_slots_6_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fp_val = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_fp_val :
    issue_slots_6_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fp_single = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_fp_single :
    issue_slots_6_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_pf_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_pf_if :
    issue_slots_6_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_ae_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_ae_if :
    issue_slots_6_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_ma_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_ma_if :
    issue_slots_6_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bp_debug_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_bp_debug_if :
    issue_slots_6_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bp_xcpt_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_bp_xcpt_if :
    issue_slots_6_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_fsrc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_fsrc :
    issue_slots_6_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_tsrc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_tsrc :
    issue_slots_6_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_clock = clock;
  assign slots_6_reset = reset;
  assign slots_6_io_grant = issue_slots_6_request & ~_T_605 & _T_608 & ~_T_587 | _T_605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_6_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_6_io_clear = _GEN_21[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_6_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_6_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_6_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_6_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_6_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_6_io_in_uop_valid = _GEN_25[1:0] == 2'h2 ? issue_slots_8_will_be_valid : _GEN_1228; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_6_io_in_uop_bits_switch = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_switch :
    issue_slots_7_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_switch_off = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_switch_off :
    issue_slots_7_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_unicore = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_unicore :
    issue_slots_7_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_shift = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_shift : issue_slots_7_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs3_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs3_rtype :
    issue_slots_7_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rflag = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_rflag : issue_slots_7_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_wflag = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_wflag : issue_slots_7_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prflag = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prflag :
    issue_slots_7_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pwflag = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_pwflag :
    issue_slots_7_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pflag_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_pflag_busy :
    issue_slots_7_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stale_pflag = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_stale_pflag :
    issue_slots_7_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_op1_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_op1_sel :
    issue_slots_7_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_op2_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_op2_sel :
    issue_slots_7_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_split_num = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_split_num :
    issue_slots_7_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_self_index = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_self_index :
    issue_slots_7_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rob_inst_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_rob_inst_idx :
    issue_slots_7_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_address_num = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_address_num :
    issue_slots_7_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uopc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_uopc : issue_slots_7_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_inst : issue_slots_7_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_inst :
    issue_slots_7_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_rvc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_rvc :
    issue_slots_7_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_pc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_pc :
    issue_slots_7_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iq_type = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iq_type :
    issue_slots_7_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fu_code = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_fu_code :
    issue_slots_7_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_br_type = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_br_type :
    issue_slots_7_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op1_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op1_sel :
    issue_slots_7_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op2_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op2_sel :
    issue_slots_7_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_imm_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_imm_sel :
    issue_slots_7_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op_fcn = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op_fcn :
    issue_slots_7_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_fcn_dw = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_fcn_dw :
    issue_slots_7_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_csr_cmd = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_csr_cmd :
    issue_slots_7_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_load = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_load :
    issue_slots_7_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_sta = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_sta :
    issue_slots_7_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_std = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_std :
    issue_slots_7_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op3_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op3_sel :
    issue_slots_7_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_state = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_state :
    issue_slots_7_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_p1_poisoned = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_p1_poisoned :
    issue_slots_7_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_p2_poisoned = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_p2_poisoned :
    issue_slots_7_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_br = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_br : issue_slots_7_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_jalr = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_jalr :
    issue_slots_7_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_jal = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_jal :
    issue_slots_7_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_sfb = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_sfb :
    issue_slots_7_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_br_mask = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_br_mask :
    issue_slots_7_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_br_tag = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_br_tag :
    issue_slots_7_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ftq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ftq_idx :
    issue_slots_7_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_edge_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_edge_inst :
    issue_slots_7_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pc_lob = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_pc_lob :
    issue_slots_7_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_taken = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_taken : issue_slots_7_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_imm_packed = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_imm_packed :
    issue_slots_7_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_csr_addr = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_csr_addr :
    issue_slots_7_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rob_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_rob_idx :
    issue_slots_7_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldq_idx :
    issue_slots_7_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_stq_idx :
    issue_slots_7_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rxq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_rxq_idx :
    issue_slots_7_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pdst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_pdst : issue_slots_7_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs1 : issue_slots_7_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs2 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs2 : issue_slots_7_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs3 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs3 : issue_slots_7_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ppred = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ppred : issue_slots_7_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs1_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs1_busy :
    issue_slots_7_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs2_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs2_busy :
    issue_slots_7_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs3_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs3_busy :
    issue_slots_7_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ppred_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ppred_busy :
    issue_slots_7_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stale_pdst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_stale_pdst :
    issue_slots_7_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_exception = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_exception :
    issue_slots_7_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_exc_cause = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_exc_cause :
    issue_slots_7_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bypassable = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_bypassable :
    issue_slots_7_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_cmd = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_cmd :
    issue_slots_7_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_size = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_size :
    issue_slots_7_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_signed = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_signed :
    issue_slots_7_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_fence = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_fence :
    issue_slots_7_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_fencei = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_fencei :
    issue_slots_7_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_amo = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_amo :
    issue_slots_7_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uses_ldq = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_uses_ldq :
    issue_slots_7_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uses_stq = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_uses_stq :
    issue_slots_7_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_sys_pc2epc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_sys_pc2epc :
    issue_slots_7_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_unique = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_unique :
    issue_slots_7_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_flush_on_commit = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_flush_on_commit :
    issue_slots_7_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst_is_rs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst_is_rs1 :
    issue_slots_7_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst : issue_slots_7_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs1 : issue_slots_7_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs2 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs2 : issue_slots_7_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs3 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs3 : issue_slots_7_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst_val = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst_val :
    issue_slots_7_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_dst_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_dst_rtype :
    issue_slots_7_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs1_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs1_rtype :
    issue_slots_7_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs2_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs2_rtype :
    issue_slots_7_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_frs3_en = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_frs3_en :
    issue_slots_7_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fp_val = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_fp_val :
    issue_slots_7_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fp_single = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_fp_single :
    issue_slots_7_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_pf_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_pf_if :
    issue_slots_7_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_ae_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_ae_if :
    issue_slots_7_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_ma_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_ma_if :
    issue_slots_7_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bp_debug_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_bp_debug_if :
    issue_slots_7_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bp_xcpt_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_bp_xcpt_if :
    issue_slots_7_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_fsrc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_fsrc :
    issue_slots_7_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_tsrc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_tsrc :
    issue_slots_7_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_clock = clock;
  assign slots_7_reset = reset;
  assign slots_7_io_grant = _T_646 & ~_T_617 | _T_635; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_7_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_7_io_clear = _GEN_23[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_7_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_7_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_7_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_7_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_7_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_7_io_in_uop_valid = _GEN_27[1:0] == 2'h2 ? issue_slots_9_will_be_valid : _GEN_1424; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_7_io_in_uop_bits_switch = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_switch :
    issue_slots_8_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_switch_off = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_switch_off :
    issue_slots_8_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_unicore = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_unicore :
    issue_slots_8_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_shift = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_shift : issue_slots_8_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs3_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs3_rtype :
    issue_slots_8_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rflag = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_rflag : issue_slots_8_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_wflag = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_wflag : issue_slots_8_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prflag = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prflag :
    issue_slots_8_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pwflag = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_pwflag :
    issue_slots_8_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pflag_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_pflag_busy :
    issue_slots_8_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stale_pflag = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_stale_pflag :
    issue_slots_8_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_op1_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_op1_sel :
    issue_slots_8_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_op2_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_op2_sel :
    issue_slots_8_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_split_num = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_split_num :
    issue_slots_8_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_self_index = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_self_index :
    issue_slots_8_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rob_inst_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_rob_inst_idx :
    issue_slots_8_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_address_num = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_address_num :
    issue_slots_8_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uopc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_uopc : issue_slots_8_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_inst : issue_slots_8_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_inst :
    issue_slots_8_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_rvc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_rvc :
    issue_slots_8_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_pc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_pc :
    issue_slots_8_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iq_type = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iq_type :
    issue_slots_8_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fu_code = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_fu_code :
    issue_slots_8_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_br_type = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_br_type :
    issue_slots_8_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op1_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op1_sel :
    issue_slots_8_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op2_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op2_sel :
    issue_slots_8_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_imm_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_imm_sel :
    issue_slots_8_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op_fcn = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op_fcn :
    issue_slots_8_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_fcn_dw = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_fcn_dw :
    issue_slots_8_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_csr_cmd = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_csr_cmd :
    issue_slots_8_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_load = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_load :
    issue_slots_8_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_sta = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_sta :
    issue_slots_8_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_std = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_std :
    issue_slots_8_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op3_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op3_sel :
    issue_slots_8_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_state = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_state :
    issue_slots_8_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_p1_poisoned = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_p1_poisoned :
    issue_slots_8_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_p2_poisoned = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_p2_poisoned :
    issue_slots_8_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_br = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_br : issue_slots_8_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_jalr = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_jalr :
    issue_slots_8_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_jal = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_jal :
    issue_slots_8_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_sfb = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_sfb :
    issue_slots_8_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_br_mask = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_br_mask :
    issue_slots_8_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_br_tag = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_br_tag :
    issue_slots_8_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ftq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ftq_idx :
    issue_slots_8_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_edge_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_edge_inst :
    issue_slots_8_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pc_lob = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_pc_lob :
    issue_slots_8_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_taken = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_taken : issue_slots_8_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_imm_packed = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_imm_packed :
    issue_slots_8_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_csr_addr = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_csr_addr :
    issue_slots_8_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rob_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_rob_idx :
    issue_slots_8_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldq_idx :
    issue_slots_8_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_stq_idx :
    issue_slots_8_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rxq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_rxq_idx :
    issue_slots_8_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pdst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_pdst : issue_slots_8_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs1 : issue_slots_8_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs2 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs2 : issue_slots_8_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs3 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs3 : issue_slots_8_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ppred = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ppred : issue_slots_8_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs1_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs1_busy :
    issue_slots_8_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs2_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs2_busy :
    issue_slots_8_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs3_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs3_busy :
    issue_slots_8_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ppred_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ppred_busy :
    issue_slots_8_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stale_pdst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_stale_pdst :
    issue_slots_8_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_exception = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_exception :
    issue_slots_8_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_exc_cause = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_exc_cause :
    issue_slots_8_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bypassable = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_bypassable :
    issue_slots_8_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_cmd = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_cmd :
    issue_slots_8_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_size = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_size :
    issue_slots_8_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_signed = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_signed :
    issue_slots_8_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_fence = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_fence :
    issue_slots_8_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_fencei = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_fencei :
    issue_slots_8_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_amo = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_amo :
    issue_slots_8_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uses_ldq = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_uses_ldq :
    issue_slots_8_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uses_stq = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_uses_stq :
    issue_slots_8_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_sys_pc2epc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_sys_pc2epc :
    issue_slots_8_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_unique = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_unique :
    issue_slots_8_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_flush_on_commit = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_flush_on_commit :
    issue_slots_8_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst_is_rs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst_is_rs1 :
    issue_slots_8_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst : issue_slots_8_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs1 : issue_slots_8_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs2 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs2 : issue_slots_8_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs3 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs3 : issue_slots_8_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst_val = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst_val :
    issue_slots_8_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_dst_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_dst_rtype :
    issue_slots_8_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs1_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs1_rtype :
    issue_slots_8_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs2_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs2_rtype :
    issue_slots_8_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_frs3_en = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_frs3_en :
    issue_slots_8_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fp_val = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_fp_val :
    issue_slots_8_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fp_single = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_fp_single :
    issue_slots_8_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_pf_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_pf_if :
    issue_slots_8_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_ae_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_ae_if :
    issue_slots_8_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_ma_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_ma_if :
    issue_slots_8_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bp_debug_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_bp_debug_if :
    issue_slots_8_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bp_xcpt_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_bp_xcpt_if :
    issue_slots_8_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_fsrc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_fsrc :
    issue_slots_8_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_tsrc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_tsrc :
    issue_slots_8_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_clock = clock;
  assign slots_8_reset = reset;
  assign slots_8_io_grant = issue_slots_8_request & ~_T_665 & _T_668 & ~_T_647 | _T_665; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_8_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_8_io_clear = _GEN_25[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_8_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_8_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_8_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_8_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_8_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_8_io_in_uop_valid = _GEN_29[1:0] == 2'h2 ? issue_slots_10_will_be_valid : _GEN_1620; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_8_io_in_uop_bits_switch = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_switch :
    issue_slots_9_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_switch_off = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_switch_off :
    issue_slots_9_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_unicore = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_unicore :
    issue_slots_9_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_shift = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_shift :
    issue_slots_9_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs3_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs3_rtype :
    issue_slots_9_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rflag = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_rflag :
    issue_slots_9_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_wflag = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_wflag :
    issue_slots_9_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prflag = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prflag :
    issue_slots_9_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pwflag = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_pwflag :
    issue_slots_9_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pflag_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_pflag_busy :
    issue_slots_9_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stale_pflag = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_stale_pflag :
    issue_slots_9_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_op1_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_op1_sel :
    issue_slots_9_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_op2_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_op2_sel :
    issue_slots_9_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_split_num = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_split_num :
    issue_slots_9_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_self_index = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_self_index :
    issue_slots_9_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rob_inst_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_rob_inst_idx :
    issue_slots_9_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_address_num = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_address_num :
    issue_slots_9_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uopc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_uopc : issue_slots_9_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_inst : issue_slots_9_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_inst :
    issue_slots_9_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_rvc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_rvc :
    issue_slots_9_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_pc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_pc :
    issue_slots_9_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iq_type = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iq_type :
    issue_slots_9_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fu_code = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_fu_code :
    issue_slots_9_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_br_type = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_br_type :
    issue_slots_9_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op1_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op1_sel :
    issue_slots_9_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op2_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op2_sel :
    issue_slots_9_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_imm_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_imm_sel :
    issue_slots_9_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op_fcn = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op_fcn :
    issue_slots_9_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_fcn_dw = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_fcn_dw :
    issue_slots_9_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_csr_cmd = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_csr_cmd :
    issue_slots_9_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_load = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_load :
    issue_slots_9_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_sta = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_sta :
    issue_slots_9_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_std = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_std :
    issue_slots_9_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op3_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op3_sel :
    issue_slots_9_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_state = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_state :
    issue_slots_9_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_p1_poisoned = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_p1_poisoned :
    issue_slots_9_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_p2_poisoned = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_p2_poisoned :
    issue_slots_9_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_br = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_br :
    issue_slots_9_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_jalr = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_jalr :
    issue_slots_9_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_jal = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_jal :
    issue_slots_9_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_sfb = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_sfb :
    issue_slots_9_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_br_mask = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_br_mask :
    issue_slots_9_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_br_tag = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_br_tag :
    issue_slots_9_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ftq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ftq_idx :
    issue_slots_9_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_edge_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_edge_inst :
    issue_slots_9_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pc_lob = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_pc_lob :
    issue_slots_9_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_taken = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_taken :
    issue_slots_9_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_imm_packed = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_imm_packed :
    issue_slots_9_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_csr_addr = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_csr_addr :
    issue_slots_9_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rob_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_rob_idx :
    issue_slots_9_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldq_idx :
    issue_slots_9_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_stq_idx :
    issue_slots_9_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rxq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_rxq_idx :
    issue_slots_9_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pdst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_pdst : issue_slots_9_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs1 : issue_slots_9_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs2 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs2 : issue_slots_9_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs3 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs3 : issue_slots_9_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ppred = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ppred :
    issue_slots_9_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs1_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs1_busy :
    issue_slots_9_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs2_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs2_busy :
    issue_slots_9_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs3_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs3_busy :
    issue_slots_9_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ppred_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ppred_busy :
    issue_slots_9_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stale_pdst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_stale_pdst :
    issue_slots_9_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_exception = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_exception :
    issue_slots_9_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_exc_cause = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_exc_cause :
    issue_slots_9_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bypassable = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_bypassable :
    issue_slots_9_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_cmd = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_cmd :
    issue_slots_9_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_size = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_size :
    issue_slots_9_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_signed = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_signed :
    issue_slots_9_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_fence = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_fence :
    issue_slots_9_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_fencei = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_fencei :
    issue_slots_9_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_amo = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_amo :
    issue_slots_9_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uses_ldq = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_uses_ldq :
    issue_slots_9_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uses_stq = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_uses_stq :
    issue_slots_9_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_sys_pc2epc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_sys_pc2epc :
    issue_slots_9_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_unique = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_unique :
    issue_slots_9_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_flush_on_commit = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_flush_on_commit :
    issue_slots_9_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst_is_rs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst_is_rs1 :
    issue_slots_9_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst : issue_slots_9_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs1 : issue_slots_9_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs2 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs2 : issue_slots_9_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs3 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs3 : issue_slots_9_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst_val = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst_val :
    issue_slots_9_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_dst_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_dst_rtype :
    issue_slots_9_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs1_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs1_rtype :
    issue_slots_9_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs2_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs2_rtype :
    issue_slots_9_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_frs3_en = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_frs3_en :
    issue_slots_9_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fp_val = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_fp_val :
    issue_slots_9_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fp_single = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_fp_single :
    issue_slots_9_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_pf_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_pf_if :
    issue_slots_9_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_ae_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_ae_if :
    issue_slots_9_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_ma_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_ma_if :
    issue_slots_9_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bp_debug_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_bp_debug_if :
    issue_slots_9_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bp_xcpt_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_bp_xcpt_if :
    issue_slots_9_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_fsrc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_fsrc :
    issue_slots_9_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_tsrc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_tsrc :
    issue_slots_9_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_clock = clock;
  assign slots_9_reset = reset;
  assign slots_9_io_grant = issue_slots_9_request & ~_T_695 & _T_698 & ~_T_677 | _T_695; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_9_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_9_io_clear = _GEN_27[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_9_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_9_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_9_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_9_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_9_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_9_io_in_uop_valid = _GEN_31[1:0] == 2'h2 ? issue_slots_11_will_be_valid : _GEN_1816; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_9_io_in_uop_bits_switch = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_switch :
    issue_slots_10_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_switch_off = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_switch_off :
    issue_slots_10_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_unicore = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_unicore :
    issue_slots_10_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_shift = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_shift :
    issue_slots_10_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs3_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs3_rtype :
    issue_slots_10_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rflag = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_rflag :
    issue_slots_10_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_wflag = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_wflag :
    issue_slots_10_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prflag = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prflag :
    issue_slots_10_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pwflag = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_pwflag :
    issue_slots_10_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pflag_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_pflag_busy :
    issue_slots_10_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stale_pflag = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_stale_pflag :
    issue_slots_10_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_op1_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_op1_sel :
    issue_slots_10_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_op2_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_op2_sel :
    issue_slots_10_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_split_num = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_split_num :
    issue_slots_10_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_self_index = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_self_index :
    issue_slots_10_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rob_inst_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_rob_inst_idx :
    issue_slots_10_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_address_num = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_address_num :
    issue_slots_10_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uopc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_uopc : issue_slots_10_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_inst : issue_slots_10_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_inst :
    issue_slots_10_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_rvc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_rvc :
    issue_slots_10_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_pc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_pc :
    issue_slots_10_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iq_type = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iq_type :
    issue_slots_10_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fu_code = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_fu_code :
    issue_slots_10_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_br_type = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_br_type :
    issue_slots_10_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op1_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op1_sel :
    issue_slots_10_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op2_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op2_sel :
    issue_slots_10_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_imm_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_imm_sel :
    issue_slots_10_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op_fcn = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op_fcn :
    issue_slots_10_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_fcn_dw = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_fcn_dw :
    issue_slots_10_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_csr_cmd = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_csr_cmd :
    issue_slots_10_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_load = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_load :
    issue_slots_10_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_sta = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_sta :
    issue_slots_10_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_std = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_std :
    issue_slots_10_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op3_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op3_sel :
    issue_slots_10_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_state = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_state :
    issue_slots_10_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_p1_poisoned = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_p1_poisoned :
    issue_slots_10_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_p2_poisoned = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_p2_poisoned :
    issue_slots_10_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_br = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_br :
    issue_slots_10_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_jalr = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_jalr :
    issue_slots_10_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_jal = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_jal :
    issue_slots_10_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_sfb = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_sfb :
    issue_slots_10_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_br_mask = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_br_mask :
    issue_slots_10_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_br_tag = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_br_tag :
    issue_slots_10_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ftq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ftq_idx :
    issue_slots_10_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_edge_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_edge_inst :
    issue_slots_10_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pc_lob = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_pc_lob :
    issue_slots_10_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_taken = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_taken :
    issue_slots_10_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_imm_packed = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_imm_packed :
    issue_slots_10_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_csr_addr = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_csr_addr :
    issue_slots_10_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rob_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_rob_idx :
    issue_slots_10_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldq_idx :
    issue_slots_10_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_stq_idx :
    issue_slots_10_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rxq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_rxq_idx :
    issue_slots_10_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pdst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_pdst : issue_slots_10_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs1 : issue_slots_10_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs2 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs2 : issue_slots_10_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs3 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs3 : issue_slots_10_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ppred = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ppred :
    issue_slots_10_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs1_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs1_busy :
    issue_slots_10_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs2_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs2_busy :
    issue_slots_10_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs3_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs3_busy :
    issue_slots_10_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ppred_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ppred_busy :
    issue_slots_10_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stale_pdst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_stale_pdst :
    issue_slots_10_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_exception = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_exception :
    issue_slots_10_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_exc_cause = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_exc_cause :
    issue_slots_10_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bypassable = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_bypassable :
    issue_slots_10_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_cmd = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_cmd :
    issue_slots_10_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_size = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_size :
    issue_slots_10_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_signed = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_signed :
    issue_slots_10_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_fence = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_fence :
    issue_slots_10_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_fencei = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_fencei :
    issue_slots_10_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_amo = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_amo :
    issue_slots_10_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uses_ldq = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_uses_ldq :
    issue_slots_10_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uses_stq = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_uses_stq :
    issue_slots_10_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_sys_pc2epc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_sys_pc2epc :
    issue_slots_10_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_unique = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_unique :
    issue_slots_10_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_flush_on_commit = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_flush_on_commit :
    issue_slots_10_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst_is_rs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst_is_rs1 :
    issue_slots_10_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst : issue_slots_10_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs1 : issue_slots_10_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs2 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs2 : issue_slots_10_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs3 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs3 : issue_slots_10_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst_val = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst_val :
    issue_slots_10_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_dst_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_dst_rtype :
    issue_slots_10_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs1_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs1_rtype :
    issue_slots_10_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs2_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs2_rtype :
    issue_slots_10_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_frs3_en = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_frs3_en :
    issue_slots_10_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fp_val = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_fp_val :
    issue_slots_10_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fp_single = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_fp_single :
    issue_slots_10_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_pf_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_pf_if :
    issue_slots_10_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_ae_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_ae_if :
    issue_slots_10_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_ma_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_ma_if :
    issue_slots_10_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bp_debug_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_bp_debug_if :
    issue_slots_10_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bp_xcpt_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_bp_xcpt_if :
    issue_slots_10_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_fsrc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_fsrc :
    issue_slots_10_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_tsrc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_tsrc :
    issue_slots_10_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_clock = clock;
  assign slots_10_reset = reset;
  assign slots_10_io_grant = issue_slots_10_request & ~_T_725 & _T_728 & ~_T_707 | _T_725; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_10_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_10_io_clear = _GEN_29[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_10_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_10_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_10_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_10_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_10_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_10_io_in_uop_valid = _GEN_33[1:0] == 2'h2 ? issue_slots_12_will_be_valid : _GEN_2012; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_10_io_in_uop_bits_switch = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_switch :
    issue_slots_11_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_switch_off = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_switch_off :
    issue_slots_11_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_unicore = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_unicore :
    issue_slots_11_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_shift = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_shift :
    issue_slots_11_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs3_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs3_rtype :
    issue_slots_11_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rflag = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_rflag :
    issue_slots_11_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_wflag = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_wflag :
    issue_slots_11_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prflag = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_prflag :
    issue_slots_11_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pwflag = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_pwflag :
    issue_slots_11_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pflag_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_pflag_busy :
    issue_slots_11_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stale_pflag = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_stale_pflag :
    issue_slots_11_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_op1_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_op1_sel :
    issue_slots_11_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_op2_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_op2_sel :
    issue_slots_11_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_split_num = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_split_num :
    issue_slots_11_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_self_index = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_self_index :
    issue_slots_11_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rob_inst_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_rob_inst_idx :
    issue_slots_11_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_address_num = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_address_num :
    issue_slots_11_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uopc = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_uopc : issue_slots_11_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_inst = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_inst : issue_slots_11_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_inst = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_inst :
    issue_slots_11_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_rvc = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_rvc :
    issue_slots_11_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_pc = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_pc :
    issue_slots_11_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iq_type = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_iq_type :
    issue_slots_11_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fu_code = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_fu_code :
    issue_slots_11_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_br_type = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_br_type :
    issue_slots_11_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op1_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op1_sel :
    issue_slots_11_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op2_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op2_sel :
    issue_slots_11_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_imm_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_imm_sel :
    issue_slots_11_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op_fcn = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op_fcn :
    issue_slots_11_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_fcn_dw = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_fcn_dw :
    issue_slots_11_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_csr_cmd = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_csr_cmd :
    issue_slots_11_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_load = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_is_load :
    issue_slots_11_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_sta = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_is_sta :
    issue_slots_11_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_std = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_is_std :
    issue_slots_11_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op3_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op3_sel :
    issue_slots_11_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_state = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_iw_state :
    issue_slots_11_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_p1_poisoned = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_iw_p1_poisoned :
    issue_slots_11_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_p2_poisoned = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_iw_p2_poisoned :
    issue_slots_11_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_br = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_br :
    issue_slots_11_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_jalr = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_jalr :
    issue_slots_11_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_jal = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_jal :
    issue_slots_11_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_sfb = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_sfb :
    issue_slots_11_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_br_mask = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_br_mask :
    issue_slots_11_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_br_tag = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_br_tag :
    issue_slots_11_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ftq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ftq_idx :
    issue_slots_11_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_edge_inst = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_edge_inst :
    issue_slots_11_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pc_lob = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_pc_lob :
    issue_slots_11_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_taken = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_taken :
    issue_slots_11_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_imm_packed = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_imm_packed :
    issue_slots_11_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_csr_addr = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_csr_addr :
    issue_slots_11_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rob_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_rob_idx :
    issue_slots_11_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ldq_idx :
    issue_slots_11_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_stq_idx :
    issue_slots_11_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rxq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_rxq_idx :
    issue_slots_11_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pdst = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_pdst : issue_slots_11_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs1 = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_prs1 : issue_slots_11_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs2 = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_prs2 : issue_slots_11_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs3 = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_prs3 : issue_slots_11_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ppred = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ppred :
    issue_slots_11_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs1_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_prs1_busy :
    issue_slots_11_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs2_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_prs2_busy :
    issue_slots_11_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs3_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_prs3_busy :
    issue_slots_11_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ppred_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ppred_busy :
    issue_slots_11_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stale_pdst = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_stale_pdst :
    issue_slots_11_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_exception = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_exception :
    issue_slots_11_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_exc_cause = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_exc_cause :
    issue_slots_11_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bypassable = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_bypassable :
    issue_slots_11_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_cmd = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_mem_cmd :
    issue_slots_11_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_size = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_mem_size :
    issue_slots_11_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_signed = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_mem_signed :
    issue_slots_11_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_fence = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_fence :
    issue_slots_11_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_fencei = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_fencei :
    issue_slots_11_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_amo = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_amo :
    issue_slots_11_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uses_ldq = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_uses_ldq :
    issue_slots_11_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uses_stq = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_uses_stq :
    issue_slots_11_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_sys_pc2epc = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_sys_pc2epc :
    issue_slots_11_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_unique = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_is_unique :
    issue_slots_11_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_flush_on_commit = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_flush_on_commit :
    issue_slots_11_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst_is_rs1 = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ldst_is_rs1 :
    issue_slots_11_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ldst : issue_slots_11_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs1 = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs1 : issue_slots_11_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs2 = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs2 : issue_slots_11_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs3 = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs3 : issue_slots_11_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst_val = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_ldst_val :
    issue_slots_11_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_dst_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_dst_rtype :
    issue_slots_11_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs1_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs1_rtype :
    issue_slots_11_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs2_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs2_rtype :
    issue_slots_11_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_frs3_en = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_frs3_en :
    issue_slots_11_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fp_val = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_fp_val :
    issue_slots_11_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fp_single = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_fp_single :
    issue_slots_11_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_pf_if = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_xcpt_pf_if :
    issue_slots_11_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_ae_if = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_xcpt_ae_if :
    issue_slots_11_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_ma_if = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_xcpt_ma_if :
    issue_slots_11_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bp_debug_if = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_bp_debug_if :
    issue_slots_11_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bp_xcpt_if = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_bp_xcpt_if :
    issue_slots_11_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_fsrc = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_fsrc :
    issue_slots_11_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_tsrc = _GEN_33[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_tsrc :
    issue_slots_11_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_clock = clock;
  assign slots_11_reset = reset;
  assign slots_11_io_grant = issue_slots_11_request & ~_T_755 & _T_758 & ~_T_737 | _T_755; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_11_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_11_io_clear = _GEN_31[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_11_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_11_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_11_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_11_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_11_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_11_io_in_uop_valid = _GEN_35[1:0] == 2'h2 ? issue_slots_13_will_be_valid : _GEN_2208; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_11_io_in_uop_bits_switch = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_switch :
    issue_slots_12_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_switch_off = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_switch_off :
    issue_slots_12_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_unicore = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_unicore :
    issue_slots_12_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_shift = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_shift :
    issue_slots_12_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs3_rtype = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs3_rtype :
    issue_slots_12_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rflag = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_rflag :
    issue_slots_12_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_wflag = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_wflag :
    issue_slots_12_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prflag = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_prflag :
    issue_slots_12_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pwflag = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_pwflag :
    issue_slots_12_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pflag_busy = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_pflag_busy :
    issue_slots_12_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stale_pflag = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_stale_pflag :
    issue_slots_12_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_op1_sel = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_op1_sel :
    issue_slots_12_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_op2_sel = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_op2_sel :
    issue_slots_12_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_split_num = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_split_num :
    issue_slots_12_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_self_index = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_self_index :
    issue_slots_12_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rob_inst_idx = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_rob_inst_idx :
    issue_slots_12_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_address_num = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_address_num :
    issue_slots_12_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uopc = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_uopc : issue_slots_12_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_inst = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_inst : issue_slots_12_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_inst = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_inst :
    issue_slots_12_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_rvc = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_rvc :
    issue_slots_12_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_pc = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_pc :
    issue_slots_12_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iq_type = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_iq_type :
    issue_slots_12_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fu_code = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_fu_code :
    issue_slots_12_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_br_type = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_br_type :
    issue_slots_12_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op1_sel = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op1_sel :
    issue_slots_12_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op2_sel = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op2_sel :
    issue_slots_12_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_imm_sel = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_imm_sel :
    issue_slots_12_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op_fcn = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op_fcn :
    issue_slots_12_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_fcn_dw = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_fcn_dw :
    issue_slots_12_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_csr_cmd = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_csr_cmd :
    issue_slots_12_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_load = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_is_load :
    issue_slots_12_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_sta = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_is_sta :
    issue_slots_12_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_std = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_is_std :
    issue_slots_12_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op3_sel = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op3_sel :
    issue_slots_12_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_state = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_iw_state :
    issue_slots_12_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_p1_poisoned = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_iw_p1_poisoned :
    issue_slots_12_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_p2_poisoned = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_iw_p2_poisoned :
    issue_slots_12_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_br = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_br :
    issue_slots_12_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_jalr = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_jalr :
    issue_slots_12_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_jal = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_jal :
    issue_slots_12_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_sfb = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_sfb :
    issue_slots_12_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_br_mask = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_br_mask :
    issue_slots_12_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_br_tag = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_br_tag :
    issue_slots_12_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ftq_idx = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ftq_idx :
    issue_slots_12_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_edge_inst = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_edge_inst :
    issue_slots_12_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pc_lob = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_pc_lob :
    issue_slots_12_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_taken = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_taken :
    issue_slots_12_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_imm_packed = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_imm_packed :
    issue_slots_12_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_csr_addr = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_csr_addr :
    issue_slots_12_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rob_idx = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_rob_idx :
    issue_slots_12_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldq_idx = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ldq_idx :
    issue_slots_12_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stq_idx = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_stq_idx :
    issue_slots_12_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rxq_idx = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_rxq_idx :
    issue_slots_12_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pdst = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_pdst : issue_slots_12_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs1 = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_prs1 : issue_slots_12_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs2 = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_prs2 : issue_slots_12_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs3 = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_prs3 : issue_slots_12_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ppred = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ppred :
    issue_slots_12_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs1_busy = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_prs1_busy :
    issue_slots_12_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs2_busy = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_prs2_busy :
    issue_slots_12_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs3_busy = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_prs3_busy :
    issue_slots_12_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ppred_busy = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ppred_busy :
    issue_slots_12_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stale_pdst = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_stale_pdst :
    issue_slots_12_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_exception = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_exception :
    issue_slots_12_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_exc_cause = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_exc_cause :
    issue_slots_12_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bypassable = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_bypassable :
    issue_slots_12_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_cmd = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_mem_cmd :
    issue_slots_12_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_size = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_mem_size :
    issue_slots_12_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_signed = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_mem_signed :
    issue_slots_12_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_fence = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_fence :
    issue_slots_12_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_fencei = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_fencei :
    issue_slots_12_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_amo = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_amo :
    issue_slots_12_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uses_ldq = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_uses_ldq :
    issue_slots_12_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uses_stq = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_uses_stq :
    issue_slots_12_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_sys_pc2epc = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_sys_pc2epc :
    issue_slots_12_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_unique = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_is_unique :
    issue_slots_12_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_flush_on_commit = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_flush_on_commit :
    issue_slots_12_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst_is_rs1 = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ldst_is_rs1 :
    issue_slots_12_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ldst : issue_slots_12_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs1 = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs1 : issue_slots_12_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs2 = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs2 : issue_slots_12_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs3 = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs3 : issue_slots_12_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst_val = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_ldst_val :
    issue_slots_12_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_dst_rtype = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_dst_rtype :
    issue_slots_12_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs1_rtype = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs1_rtype :
    issue_slots_12_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs2_rtype = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs2_rtype :
    issue_slots_12_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_frs3_en = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_frs3_en :
    issue_slots_12_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fp_val = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_fp_val :
    issue_slots_12_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fp_single = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_fp_single :
    issue_slots_12_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_pf_if = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_xcpt_pf_if :
    issue_slots_12_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_ae_if = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_xcpt_ae_if :
    issue_slots_12_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_ma_if = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_xcpt_ma_if :
    issue_slots_12_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bp_debug_if = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_bp_debug_if :
    issue_slots_12_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bp_xcpt_if = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_bp_xcpt_if :
    issue_slots_12_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_fsrc = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_fsrc :
    issue_slots_12_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_tsrc = _GEN_35[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_tsrc :
    issue_slots_12_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_clock = clock;
  assign slots_12_reset = reset;
  assign slots_12_io_grant = _T_796 & ~_T_767 | _T_785; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_12_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_12_io_clear = _GEN_33[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_12_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_12_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_12_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_12_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_12_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_12_io_in_uop_valid = _GEN_37[1:0] == 2'h2 ? issue_slots_14_will_be_valid : _GEN_2404; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_12_io_in_uop_bits_switch = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_switch :
    issue_slots_13_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_switch_off = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_switch_off :
    issue_slots_13_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_unicore = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_unicore :
    issue_slots_13_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_shift = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_shift :
    issue_slots_13_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs3_rtype = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs3_rtype :
    issue_slots_13_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rflag = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_rflag :
    issue_slots_13_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_wflag = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_wflag :
    issue_slots_13_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prflag = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_prflag :
    issue_slots_13_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pwflag = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_pwflag :
    issue_slots_13_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pflag_busy = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_pflag_busy :
    issue_slots_13_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_stale_pflag = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_stale_pflag :
    issue_slots_13_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_op1_sel = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_op1_sel :
    issue_slots_13_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_op2_sel = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_op2_sel :
    issue_slots_13_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_split_num = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_split_num :
    issue_slots_13_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_self_index = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_self_index :
    issue_slots_13_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rob_inst_idx = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_rob_inst_idx :
    issue_slots_13_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_address_num = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_address_num :
    issue_slots_13_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_uopc = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_uopc : issue_slots_13_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_inst = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_inst : issue_slots_13_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_inst = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_inst :
    issue_slots_13_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_rvc = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_rvc :
    issue_slots_13_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_pc = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_pc :
    issue_slots_13_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iq_type = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_iq_type :
    issue_slots_13_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_fu_code = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_fu_code :
    issue_slots_13_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_br_type = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_br_type :
    issue_slots_13_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op1_sel = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op1_sel :
    issue_slots_13_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op2_sel = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op2_sel :
    issue_slots_13_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_imm_sel = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_imm_sel :
    issue_slots_13_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op_fcn = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op_fcn :
    issue_slots_13_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_fcn_dw = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_fcn_dw :
    issue_slots_13_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_csr_cmd = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_csr_cmd :
    issue_slots_13_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_is_load = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_is_load :
    issue_slots_13_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_is_sta = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_is_sta :
    issue_slots_13_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_is_std = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_is_std :
    issue_slots_13_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op3_sel = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op3_sel :
    issue_slots_13_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iw_state = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_iw_state :
    issue_slots_13_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iw_p1_poisoned = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_iw_p1_poisoned :
    issue_slots_13_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iw_p2_poisoned = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_iw_p2_poisoned :
    issue_slots_13_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_br = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_br :
    issue_slots_13_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_jalr = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_jalr :
    issue_slots_13_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_jal = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_jal :
    issue_slots_13_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_sfb = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_sfb :
    issue_slots_13_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_br_mask = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_br_mask :
    issue_slots_13_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_br_tag = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_br_tag :
    issue_slots_13_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ftq_idx = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ftq_idx :
    issue_slots_13_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_edge_inst = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_edge_inst :
    issue_slots_13_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pc_lob = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_pc_lob :
    issue_slots_13_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_taken = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_taken :
    issue_slots_13_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_imm_packed = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_imm_packed :
    issue_slots_13_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_csr_addr = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_csr_addr :
    issue_slots_13_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rob_idx = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_rob_idx :
    issue_slots_13_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldq_idx = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ldq_idx :
    issue_slots_13_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_stq_idx = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_stq_idx :
    issue_slots_13_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rxq_idx = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_rxq_idx :
    issue_slots_13_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pdst = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_pdst : issue_slots_13_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs1 = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_prs1 : issue_slots_13_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs2 = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_prs2 : issue_slots_13_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs3 = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_prs3 : issue_slots_13_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ppred = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ppred :
    issue_slots_13_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs1_busy = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_prs1_busy :
    issue_slots_13_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs2_busy = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_prs2_busy :
    issue_slots_13_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs3_busy = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_prs3_busy :
    issue_slots_13_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ppred_busy = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ppred_busy :
    issue_slots_13_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_stale_pdst = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_stale_pdst :
    issue_slots_13_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_exception = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_exception :
    issue_slots_13_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_exc_cause = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_exc_cause :
    issue_slots_13_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_bypassable = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_bypassable :
    issue_slots_13_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_mem_cmd = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_mem_cmd :
    issue_slots_13_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_mem_size = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_mem_size :
    issue_slots_13_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_mem_signed = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_mem_signed :
    issue_slots_13_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_fence = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_fence :
    issue_slots_13_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_fencei = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_fencei :
    issue_slots_13_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_amo = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_amo :
    issue_slots_13_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_uses_ldq = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_uses_ldq :
    issue_slots_13_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_uses_stq = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_uses_stq :
    issue_slots_13_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_sys_pc2epc = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_sys_pc2epc :
    issue_slots_13_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_unique = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_is_unique :
    issue_slots_13_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_flush_on_commit = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_flush_on_commit :
    issue_slots_13_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldst_is_rs1 = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ldst_is_rs1 :
    issue_slots_13_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldst = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ldst : issue_slots_13_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs1 = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs1 : issue_slots_13_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs2 = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs2 : issue_slots_13_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs3 = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs3 : issue_slots_13_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldst_val = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_ldst_val :
    issue_slots_13_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_dst_rtype = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_dst_rtype :
    issue_slots_13_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs1_rtype = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs1_rtype :
    issue_slots_13_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs2_rtype = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs2_rtype :
    issue_slots_13_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_frs3_en = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_frs3_en :
    issue_slots_13_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_fp_val = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_fp_val :
    issue_slots_13_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_fp_single = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_fp_single :
    issue_slots_13_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_xcpt_pf_if = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_xcpt_pf_if :
    issue_slots_13_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_xcpt_ae_if = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_xcpt_ae_if :
    issue_slots_13_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_xcpt_ma_if = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_xcpt_ma_if :
    issue_slots_13_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_bp_debug_if = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_bp_debug_if :
    issue_slots_13_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_bp_xcpt_if = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_bp_xcpt_if :
    issue_slots_13_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_fsrc = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_fsrc :
    issue_slots_13_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_tsrc = _GEN_37[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_tsrc :
    issue_slots_13_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_clock = clock;
  assign slots_13_reset = reset;
  assign slots_13_io_grant = issue_slots_13_request & ~_T_815 & _T_818 & ~_T_797 | _T_815; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_13_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_13_io_clear = _GEN_35[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_13_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_13_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_13_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_13_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_13_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_13_io_in_uop_valid = _GEN_39[1:0] == 2'h2 ? issue_slots_15_will_be_valid : _GEN_2600; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_13_io_in_uop_bits_switch = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_switch :
    issue_slots_14_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_switch_off = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_switch_off :
    issue_slots_14_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_unicore = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_unicore :
    issue_slots_14_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_shift = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_shift :
    issue_slots_14_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs3_rtype = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs3_rtype :
    issue_slots_14_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rflag = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_rflag :
    issue_slots_14_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_wflag = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_wflag :
    issue_slots_14_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prflag = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_prflag :
    issue_slots_14_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pwflag = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_pwflag :
    issue_slots_14_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pflag_busy = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_pflag_busy :
    issue_slots_14_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_stale_pflag = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_stale_pflag :
    issue_slots_14_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_op1_sel = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_op1_sel :
    issue_slots_14_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_op2_sel = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_op2_sel :
    issue_slots_14_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_split_num = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_split_num :
    issue_slots_14_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_self_index = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_self_index :
    issue_slots_14_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rob_inst_idx = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_rob_inst_idx :
    issue_slots_14_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_address_num = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_address_num :
    issue_slots_14_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_uopc = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_uopc : issue_slots_14_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_inst = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_inst : issue_slots_14_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_inst = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_inst :
    issue_slots_14_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_rvc = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_rvc :
    issue_slots_14_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_pc = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_pc :
    issue_slots_14_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iq_type = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_iq_type :
    issue_slots_14_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_fu_code = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_fu_code :
    issue_slots_14_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_br_type = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_br_type :
    issue_slots_14_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op1_sel = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op1_sel :
    issue_slots_14_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op2_sel = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op2_sel :
    issue_slots_14_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_imm_sel = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_imm_sel :
    issue_slots_14_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op_fcn = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op_fcn :
    issue_slots_14_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_fcn_dw = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_fcn_dw :
    issue_slots_14_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_csr_cmd = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_csr_cmd :
    issue_slots_14_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_is_load = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_is_load :
    issue_slots_14_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_is_sta = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_is_sta :
    issue_slots_14_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_is_std = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_is_std :
    issue_slots_14_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op3_sel = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op3_sel :
    issue_slots_14_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iw_state = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_iw_state :
    issue_slots_14_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iw_p1_poisoned = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_iw_p1_poisoned :
    issue_slots_14_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iw_p2_poisoned = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_iw_p2_poisoned :
    issue_slots_14_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_br = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_br :
    issue_slots_14_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_jalr = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_jalr :
    issue_slots_14_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_jal = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_jal :
    issue_slots_14_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_sfb = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_sfb :
    issue_slots_14_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_br_mask = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_br_mask :
    issue_slots_14_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_br_tag = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_br_tag :
    issue_slots_14_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ftq_idx = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ftq_idx :
    issue_slots_14_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_edge_inst = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_edge_inst :
    issue_slots_14_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pc_lob = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_pc_lob :
    issue_slots_14_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_taken = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_taken :
    issue_slots_14_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_imm_packed = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_imm_packed :
    issue_slots_14_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_csr_addr = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_csr_addr :
    issue_slots_14_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rob_idx = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_rob_idx :
    issue_slots_14_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldq_idx = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ldq_idx :
    issue_slots_14_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_stq_idx = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_stq_idx :
    issue_slots_14_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rxq_idx = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_rxq_idx :
    issue_slots_14_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pdst = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_pdst : issue_slots_14_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs1 = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_prs1 : issue_slots_14_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs2 = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_prs2 : issue_slots_14_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs3 = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_prs3 : issue_slots_14_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ppred = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ppred :
    issue_slots_14_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs1_busy = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_prs1_busy :
    issue_slots_14_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs2_busy = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_prs2_busy :
    issue_slots_14_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs3_busy = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_prs3_busy :
    issue_slots_14_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ppred_busy = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ppred_busy :
    issue_slots_14_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_stale_pdst = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_stale_pdst :
    issue_slots_14_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_exception = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_exception :
    issue_slots_14_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_exc_cause = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_exc_cause :
    issue_slots_14_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_bypassable = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_bypassable :
    issue_slots_14_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_mem_cmd = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_mem_cmd :
    issue_slots_14_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_mem_size = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_mem_size :
    issue_slots_14_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_mem_signed = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_mem_signed :
    issue_slots_14_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_fence = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_fence :
    issue_slots_14_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_fencei = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_fencei :
    issue_slots_14_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_amo = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_amo :
    issue_slots_14_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_uses_ldq = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_uses_ldq :
    issue_slots_14_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_uses_stq = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_uses_stq :
    issue_slots_14_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_sys_pc2epc = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_sys_pc2epc :
    issue_slots_14_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_unique = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_is_unique :
    issue_slots_14_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_flush_on_commit = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_flush_on_commit :
    issue_slots_14_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldst_is_rs1 = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ldst_is_rs1 :
    issue_slots_14_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldst = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ldst : issue_slots_14_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs1 = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs1 : issue_slots_14_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs2 = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs2 : issue_slots_14_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs3 = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs3 : issue_slots_14_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldst_val = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_ldst_val :
    issue_slots_14_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_dst_rtype = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_dst_rtype :
    issue_slots_14_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs1_rtype = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs1_rtype :
    issue_slots_14_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs2_rtype = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs2_rtype :
    issue_slots_14_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_frs3_en = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_frs3_en :
    issue_slots_14_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_fp_val = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_fp_val :
    issue_slots_14_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_fp_single = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_fp_single :
    issue_slots_14_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_xcpt_pf_if = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_xcpt_pf_if :
    issue_slots_14_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_xcpt_ae_if = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_xcpt_ae_if :
    issue_slots_14_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_xcpt_ma_if = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_xcpt_ma_if :
    issue_slots_14_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_bp_debug_if = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_bp_debug_if :
    issue_slots_14_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_bp_xcpt_if = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_bp_xcpt_if :
    issue_slots_14_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_fsrc = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_fsrc :
    issue_slots_14_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_tsrc = _GEN_39[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_tsrc :
    issue_slots_14_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_clock = clock;
  assign slots_14_reset = reset;
  assign slots_14_io_grant = issue_slots_14_request & ~_T_845 & _T_848 & ~_T_827 | _T_845; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_14_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_14_io_clear = _GEN_37[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_14_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_14_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_14_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_14_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_14_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_14_io_in_uop_valid = _GEN_41[1:0] == 2'h2 ? issue_slots_16_will_be_valid : _GEN_2796; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_14_io_in_uop_bits_switch = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_switch :
    issue_slots_15_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_switch_off = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_switch_off :
    issue_slots_15_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_unicore = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_unicore :
    issue_slots_15_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_shift = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_shift :
    issue_slots_15_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs3_rtype = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_lrs3_rtype :
    issue_slots_15_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rflag = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_rflag :
    issue_slots_15_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_wflag = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_wflag :
    issue_slots_15_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prflag = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_prflag :
    issue_slots_15_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pwflag = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_pwflag :
    issue_slots_15_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pflag_busy = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_pflag_busy :
    issue_slots_15_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_stale_pflag = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_stale_pflag :
    issue_slots_15_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_op1_sel = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_op1_sel :
    issue_slots_15_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_op2_sel = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_op2_sel :
    issue_slots_15_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_split_num = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_split_num :
    issue_slots_15_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_self_index = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_self_index :
    issue_slots_15_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rob_inst_idx = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_rob_inst_idx :
    issue_slots_15_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_address_num = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_address_num :
    issue_slots_15_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_uopc = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_uopc : issue_slots_15_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_inst = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_inst : issue_slots_15_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_inst = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_debug_inst :
    issue_slots_15_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_rvc = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_rvc :
    issue_slots_15_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_pc = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_debug_pc :
    issue_slots_15_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iq_type = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_iq_type :
    issue_slots_15_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_fu_code = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_fu_code :
    issue_slots_15_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_br_type = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_br_type :
    issue_slots_15_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op1_sel = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_op1_sel :
    issue_slots_15_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op2_sel = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_op2_sel :
    issue_slots_15_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_imm_sel = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_imm_sel :
    issue_slots_15_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op_fcn = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_op_fcn :
    issue_slots_15_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_fcn_dw = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_fcn_dw :
    issue_slots_15_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_csr_cmd = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_csr_cmd :
    issue_slots_15_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_is_load = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_is_load :
    issue_slots_15_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_is_sta = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_is_sta :
    issue_slots_15_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_is_std = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_is_std :
    issue_slots_15_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op3_sel = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ctrl_op3_sel :
    issue_slots_15_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iw_state = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_iw_state :
    issue_slots_15_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iw_p1_poisoned = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_iw_p1_poisoned :
    issue_slots_15_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iw_p2_poisoned = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_iw_p2_poisoned :
    issue_slots_15_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_br = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_br :
    issue_slots_15_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_jalr = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_jalr :
    issue_slots_15_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_jal = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_jal :
    issue_slots_15_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_sfb = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_sfb :
    issue_slots_15_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_br_mask = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_br_mask :
    issue_slots_15_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_br_tag = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_br_tag :
    issue_slots_15_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ftq_idx = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ftq_idx :
    issue_slots_15_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_edge_inst = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_edge_inst :
    issue_slots_15_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pc_lob = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_pc_lob :
    issue_slots_15_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_taken = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_taken :
    issue_slots_15_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_imm_packed = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_imm_packed :
    issue_slots_15_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_csr_addr = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_csr_addr :
    issue_slots_15_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rob_idx = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_rob_idx :
    issue_slots_15_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldq_idx = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ldq_idx :
    issue_slots_15_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_stq_idx = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_stq_idx :
    issue_slots_15_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rxq_idx = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_rxq_idx :
    issue_slots_15_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pdst = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_pdst : issue_slots_15_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs1 = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_prs1 : issue_slots_15_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs2 = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_prs2 : issue_slots_15_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs3 = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_prs3 : issue_slots_15_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ppred = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ppred :
    issue_slots_15_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs1_busy = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_prs1_busy :
    issue_slots_15_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs2_busy = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_prs2_busy :
    issue_slots_15_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs3_busy = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_prs3_busy :
    issue_slots_15_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ppred_busy = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ppred_busy :
    issue_slots_15_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_stale_pdst = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_stale_pdst :
    issue_slots_15_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_exception = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_exception :
    issue_slots_15_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_exc_cause = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_exc_cause :
    issue_slots_15_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_bypassable = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_bypassable :
    issue_slots_15_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_mem_cmd = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_mem_cmd :
    issue_slots_15_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_mem_size = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_mem_size :
    issue_slots_15_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_mem_signed = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_mem_signed :
    issue_slots_15_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_fence = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_fence :
    issue_slots_15_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_fencei = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_fencei :
    issue_slots_15_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_amo = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_amo :
    issue_slots_15_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_uses_ldq = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_uses_ldq :
    issue_slots_15_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_uses_stq = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_uses_stq :
    issue_slots_15_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_sys_pc2epc = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_sys_pc2epc :
    issue_slots_15_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_unique = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_is_unique :
    issue_slots_15_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_flush_on_commit = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_flush_on_commit :
    issue_slots_15_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldst_is_rs1 = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ldst_is_rs1 :
    issue_slots_15_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldst = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ldst : issue_slots_15_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs1 = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_lrs1 : issue_slots_15_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs2 = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_lrs2 : issue_slots_15_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs3 = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_lrs3 : issue_slots_15_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldst_val = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_ldst_val :
    issue_slots_15_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_dst_rtype = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_dst_rtype :
    issue_slots_15_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs1_rtype = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_lrs1_rtype :
    issue_slots_15_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs2_rtype = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_lrs2_rtype :
    issue_slots_15_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_frs3_en = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_frs3_en :
    issue_slots_15_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_fp_val = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_fp_val :
    issue_slots_15_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_fp_single = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_fp_single :
    issue_slots_15_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_xcpt_pf_if = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_xcpt_pf_if :
    issue_slots_15_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_xcpt_ae_if = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_xcpt_ae_if :
    issue_slots_15_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_xcpt_ma_if = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_xcpt_ma_if :
    issue_slots_15_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_bp_debug_if = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_bp_debug_if :
    issue_slots_15_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_bp_xcpt_if = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_bp_xcpt_if :
    issue_slots_15_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_fsrc = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_debug_fsrc :
    issue_slots_15_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_tsrc = _GEN_41[1:0] == 2'h2 ? issue_slots_16_out_uop_debug_tsrc :
    issue_slots_15_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_clock = clock;
  assign slots_15_reset = reset;
  assign slots_15_io_grant = issue_slots_15_request & ~_T_875 & _T_878 & ~_T_857 | _T_875; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_15_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_15_io_clear = _GEN_39[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_15_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_15_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_15_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_15_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_15_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_15_io_in_uop_valid = _GEN_43[1:0] == 2'h2 ? issue_slots_17_will_be_valid : _GEN_2992; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_15_io_in_uop_bits_switch = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_switch :
    issue_slots_16_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_switch_off = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_switch_off :
    issue_slots_16_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_unicore = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_unicore :
    issue_slots_16_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_shift = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_shift :
    issue_slots_16_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs3_rtype = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_lrs3_rtype :
    issue_slots_16_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rflag = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_rflag :
    issue_slots_16_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_wflag = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_wflag :
    issue_slots_16_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prflag = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_prflag :
    issue_slots_16_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pwflag = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_pwflag :
    issue_slots_16_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pflag_busy = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_pflag_busy :
    issue_slots_16_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_stale_pflag = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_stale_pflag :
    issue_slots_16_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_op1_sel = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_op1_sel :
    issue_slots_16_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_op2_sel = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_op2_sel :
    issue_slots_16_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_split_num = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_split_num :
    issue_slots_16_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_self_index = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_self_index :
    issue_slots_16_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rob_inst_idx = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_rob_inst_idx :
    issue_slots_16_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_address_num = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_address_num :
    issue_slots_16_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_uopc = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_uopc : issue_slots_16_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_inst = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_inst : issue_slots_16_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_inst = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_debug_inst :
    issue_slots_16_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_rvc = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_rvc :
    issue_slots_16_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_pc = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_debug_pc :
    issue_slots_16_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iq_type = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_iq_type :
    issue_slots_16_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_fu_code = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_fu_code :
    issue_slots_16_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_br_type = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_br_type :
    issue_slots_16_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op1_sel = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_op1_sel :
    issue_slots_16_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op2_sel = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_op2_sel :
    issue_slots_16_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_imm_sel = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_imm_sel :
    issue_slots_16_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op_fcn = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_op_fcn :
    issue_slots_16_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_fcn_dw = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_fcn_dw :
    issue_slots_16_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_csr_cmd = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_csr_cmd :
    issue_slots_16_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_is_load = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_is_load :
    issue_slots_16_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_is_sta = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_is_sta :
    issue_slots_16_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_is_std = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_is_std :
    issue_slots_16_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op3_sel = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ctrl_op3_sel :
    issue_slots_16_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iw_state = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_iw_state :
    issue_slots_16_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iw_p1_poisoned = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_iw_p1_poisoned :
    issue_slots_16_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iw_p2_poisoned = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_iw_p2_poisoned :
    issue_slots_16_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_br = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_br :
    issue_slots_16_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_jalr = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_jalr :
    issue_slots_16_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_jal = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_jal :
    issue_slots_16_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_sfb = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_sfb :
    issue_slots_16_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_br_mask = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_br_mask :
    issue_slots_16_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_br_tag = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_br_tag :
    issue_slots_16_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ftq_idx = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ftq_idx :
    issue_slots_16_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_edge_inst = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_edge_inst :
    issue_slots_16_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pc_lob = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_pc_lob :
    issue_slots_16_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_taken = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_taken :
    issue_slots_16_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_imm_packed = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_imm_packed :
    issue_slots_16_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_csr_addr = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_csr_addr :
    issue_slots_16_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rob_idx = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_rob_idx :
    issue_slots_16_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldq_idx = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ldq_idx :
    issue_slots_16_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_stq_idx = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_stq_idx :
    issue_slots_16_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rxq_idx = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_rxq_idx :
    issue_slots_16_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pdst = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_pdst : issue_slots_16_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs1 = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_prs1 : issue_slots_16_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs2 = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_prs2 : issue_slots_16_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs3 = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_prs3 : issue_slots_16_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ppred = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ppred :
    issue_slots_16_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs1_busy = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_prs1_busy :
    issue_slots_16_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs2_busy = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_prs2_busy :
    issue_slots_16_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs3_busy = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_prs3_busy :
    issue_slots_16_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ppred_busy = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ppred_busy :
    issue_slots_16_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_stale_pdst = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_stale_pdst :
    issue_slots_16_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_exception = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_exception :
    issue_slots_16_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_exc_cause = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_exc_cause :
    issue_slots_16_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_bypassable = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_bypassable :
    issue_slots_16_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_mem_cmd = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_mem_cmd :
    issue_slots_16_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_mem_size = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_mem_size :
    issue_slots_16_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_mem_signed = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_mem_signed :
    issue_slots_16_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_fence = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_fence :
    issue_slots_16_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_fencei = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_fencei :
    issue_slots_16_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_amo = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_amo :
    issue_slots_16_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_uses_ldq = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_uses_ldq :
    issue_slots_16_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_uses_stq = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_uses_stq :
    issue_slots_16_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_sys_pc2epc = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_sys_pc2epc :
    issue_slots_16_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_unique = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_is_unique :
    issue_slots_16_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_flush_on_commit = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_flush_on_commit :
    issue_slots_16_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldst_is_rs1 = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ldst_is_rs1 :
    issue_slots_16_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldst = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ldst : issue_slots_16_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs1 = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_lrs1 : issue_slots_16_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs2 = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_lrs2 : issue_slots_16_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs3 = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_lrs3 : issue_slots_16_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldst_val = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_ldst_val :
    issue_slots_16_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_dst_rtype = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_dst_rtype :
    issue_slots_16_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs1_rtype = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_lrs1_rtype :
    issue_slots_16_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs2_rtype = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_lrs2_rtype :
    issue_slots_16_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_frs3_en = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_frs3_en :
    issue_slots_16_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_fp_val = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_fp_val :
    issue_slots_16_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_fp_single = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_fp_single :
    issue_slots_16_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_xcpt_pf_if = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_xcpt_pf_if :
    issue_slots_16_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_xcpt_ae_if = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_xcpt_ae_if :
    issue_slots_16_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_xcpt_ma_if = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_xcpt_ma_if :
    issue_slots_16_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_bp_debug_if = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_bp_debug_if :
    issue_slots_16_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_bp_xcpt_if = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_bp_xcpt_if :
    issue_slots_16_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_fsrc = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_debug_fsrc :
    issue_slots_16_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_tsrc = _GEN_43[1:0] == 2'h2 ? issue_slots_17_out_uop_debug_tsrc :
    issue_slots_16_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_clock = clock;
  assign slots_16_reset = reset;
  assign slots_16_io_grant = issue_slots_16_request & ~_T_905 & _T_908 & ~_T_887 | _T_905; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_16_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_16_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_16_io_clear = _GEN_41[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_16_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_16_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_16_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_16_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_16_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_16_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_16_io_in_uop_valid = _GEN_45[1:0] == 2'h2 ? issue_slots_18_will_be_valid : _GEN_3188; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_16_io_in_uop_bits_switch = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_switch :
    issue_slots_17_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_switch_off = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_switch_off :
    issue_slots_17_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_unicore = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_unicore :
    issue_slots_17_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_shift = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_shift :
    issue_slots_17_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_lrs3_rtype = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_lrs3_rtype :
    issue_slots_17_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_rflag = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_rflag :
    issue_slots_17_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_wflag = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_wflag :
    issue_slots_17_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_prflag = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_prflag :
    issue_slots_17_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_pwflag = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_pwflag :
    issue_slots_17_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_pflag_busy = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_pflag_busy :
    issue_slots_17_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_stale_pflag = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_stale_pflag :
    issue_slots_17_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_op1_sel = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_op1_sel :
    issue_slots_17_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_op2_sel = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_op2_sel :
    issue_slots_17_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_split_num = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_split_num :
    issue_slots_17_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_self_index = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_self_index :
    issue_slots_17_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_rob_inst_idx = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_rob_inst_idx :
    issue_slots_17_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_address_num = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_address_num :
    issue_slots_17_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_uopc = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_uopc : issue_slots_17_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_inst = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_inst : issue_slots_17_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_debug_inst = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_debug_inst :
    issue_slots_17_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_rvc = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_rvc :
    issue_slots_17_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_debug_pc = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_debug_pc :
    issue_slots_17_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_iq_type = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_iq_type :
    issue_slots_17_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_fu_code = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_fu_code :
    issue_slots_17_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_br_type = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_br_type :
    issue_slots_17_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_op1_sel = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_op1_sel :
    issue_slots_17_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_op2_sel = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_op2_sel :
    issue_slots_17_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_imm_sel = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_imm_sel :
    issue_slots_17_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_op_fcn = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_op_fcn :
    issue_slots_17_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_fcn_dw = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_fcn_dw :
    issue_slots_17_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_csr_cmd = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_csr_cmd :
    issue_slots_17_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_is_load = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_is_load :
    issue_slots_17_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_is_sta = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_is_sta :
    issue_slots_17_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_is_std = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_is_std :
    issue_slots_17_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ctrl_op3_sel = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ctrl_op3_sel :
    issue_slots_17_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_iw_state = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_iw_state :
    issue_slots_17_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_iw_p1_poisoned = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_iw_p1_poisoned :
    issue_slots_17_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_iw_p2_poisoned = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_iw_p2_poisoned :
    issue_slots_17_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_br = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_br :
    issue_slots_17_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_jalr = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_jalr :
    issue_slots_17_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_jal = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_jal :
    issue_slots_17_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_sfb = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_sfb :
    issue_slots_17_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_br_mask = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_br_mask :
    issue_slots_17_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_br_tag = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_br_tag :
    issue_slots_17_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ftq_idx = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ftq_idx :
    issue_slots_17_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_edge_inst = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_edge_inst :
    issue_slots_17_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_pc_lob = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_pc_lob :
    issue_slots_17_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_taken = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_taken :
    issue_slots_17_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_imm_packed = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_imm_packed :
    issue_slots_17_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_csr_addr = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_csr_addr :
    issue_slots_17_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_rob_idx = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_rob_idx :
    issue_slots_17_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ldq_idx = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ldq_idx :
    issue_slots_17_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_stq_idx = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_stq_idx :
    issue_slots_17_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_rxq_idx = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_rxq_idx :
    issue_slots_17_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_pdst = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_pdst : issue_slots_17_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_prs1 = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_prs1 : issue_slots_17_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_prs2 = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_prs2 : issue_slots_17_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_prs3 = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_prs3 : issue_slots_17_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ppred = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ppred :
    issue_slots_17_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_prs1_busy = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_prs1_busy :
    issue_slots_17_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_prs2_busy = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_prs2_busy :
    issue_slots_17_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_prs3_busy = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_prs3_busy :
    issue_slots_17_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ppred_busy = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ppred_busy :
    issue_slots_17_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_stale_pdst = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_stale_pdst :
    issue_slots_17_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_exception = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_exception :
    issue_slots_17_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_exc_cause = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_exc_cause :
    issue_slots_17_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_bypassable = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_bypassable :
    issue_slots_17_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_mem_cmd = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_mem_cmd :
    issue_slots_17_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_mem_size = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_mem_size :
    issue_slots_17_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_mem_signed = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_mem_signed :
    issue_slots_17_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_fence = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_fence :
    issue_slots_17_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_fencei = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_fencei :
    issue_slots_17_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_amo = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_amo :
    issue_slots_17_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_uses_ldq = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_uses_ldq :
    issue_slots_17_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_uses_stq = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_uses_stq :
    issue_slots_17_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_sys_pc2epc = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_sys_pc2epc :
    issue_slots_17_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_is_unique = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_is_unique :
    issue_slots_17_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_flush_on_commit = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_flush_on_commit :
    issue_slots_17_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ldst_is_rs1 = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ldst_is_rs1 :
    issue_slots_17_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ldst = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ldst : issue_slots_17_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_lrs1 = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_lrs1 : issue_slots_17_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_lrs2 = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_lrs2 : issue_slots_17_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_lrs3 = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_lrs3 : issue_slots_17_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_ldst_val = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_ldst_val :
    issue_slots_17_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_dst_rtype = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_dst_rtype :
    issue_slots_17_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_lrs1_rtype = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_lrs1_rtype :
    issue_slots_17_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_lrs2_rtype = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_lrs2_rtype :
    issue_slots_17_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_frs3_en = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_frs3_en :
    issue_slots_17_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_fp_val = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_fp_val :
    issue_slots_17_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_fp_single = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_fp_single :
    issue_slots_17_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_xcpt_pf_if = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_xcpt_pf_if :
    issue_slots_17_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_xcpt_ae_if = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_xcpt_ae_if :
    issue_slots_17_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_xcpt_ma_if = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_xcpt_ma_if :
    issue_slots_17_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_bp_debug_if = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_bp_debug_if :
    issue_slots_17_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_bp_xcpt_if = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_bp_xcpt_if :
    issue_slots_17_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_debug_fsrc = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_debug_fsrc :
    issue_slots_17_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_16_io_in_uop_bits_debug_tsrc = _GEN_45[1:0] == 2'h2 ? issue_slots_18_out_uop_debug_tsrc :
    issue_slots_17_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_clock = clock;
  assign slots_17_reset = reset;
  assign slots_17_io_grant = _T_946 & ~_T_917 | _T_935; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_17_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_17_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_17_io_clear = _GEN_43[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_17_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_17_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_17_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_17_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_17_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_17_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_17_io_in_uop_valid = _GEN_47[1:0] == 2'h2 ? issue_slots_19_will_be_valid : _GEN_3384; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_17_io_in_uop_bits_switch = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_switch :
    issue_slots_18_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_switch_off = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_switch_off :
    issue_slots_18_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_unicore = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_unicore :
    issue_slots_18_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_shift = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_shift :
    issue_slots_18_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_lrs3_rtype = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_lrs3_rtype :
    issue_slots_18_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_rflag = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_rflag :
    issue_slots_18_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_wflag = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_wflag :
    issue_slots_18_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_prflag = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_prflag :
    issue_slots_18_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_pwflag = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_pwflag :
    issue_slots_18_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_pflag_busy = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_pflag_busy :
    issue_slots_18_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_stale_pflag = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_stale_pflag :
    issue_slots_18_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_op1_sel = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_op1_sel :
    issue_slots_18_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_op2_sel = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_op2_sel :
    issue_slots_18_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_split_num = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_split_num :
    issue_slots_18_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_self_index = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_self_index :
    issue_slots_18_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_rob_inst_idx = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_rob_inst_idx :
    issue_slots_18_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_address_num = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_address_num :
    issue_slots_18_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_uopc = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_uopc : issue_slots_18_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_inst = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_inst : issue_slots_18_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_debug_inst = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_debug_inst :
    issue_slots_18_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_rvc = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_rvc :
    issue_slots_18_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_debug_pc = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_debug_pc :
    issue_slots_18_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_iq_type = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_iq_type :
    issue_slots_18_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_fu_code = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_fu_code :
    issue_slots_18_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_br_type = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_br_type :
    issue_slots_18_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_op1_sel = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_op1_sel :
    issue_slots_18_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_op2_sel = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_op2_sel :
    issue_slots_18_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_imm_sel = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_imm_sel :
    issue_slots_18_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_op_fcn = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_op_fcn :
    issue_slots_18_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_fcn_dw = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_fcn_dw :
    issue_slots_18_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_csr_cmd = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_csr_cmd :
    issue_slots_18_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_is_load = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_is_load :
    issue_slots_18_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_is_sta = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_is_sta :
    issue_slots_18_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_is_std = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_is_std :
    issue_slots_18_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ctrl_op3_sel = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ctrl_op3_sel :
    issue_slots_18_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_iw_state = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_iw_state :
    issue_slots_18_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_iw_p1_poisoned = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_iw_p1_poisoned :
    issue_slots_18_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_iw_p2_poisoned = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_iw_p2_poisoned :
    issue_slots_18_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_br = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_br :
    issue_slots_18_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_jalr = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_jalr :
    issue_slots_18_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_jal = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_jal :
    issue_slots_18_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_sfb = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_sfb :
    issue_slots_18_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_br_mask = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_br_mask :
    issue_slots_18_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_br_tag = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_br_tag :
    issue_slots_18_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ftq_idx = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ftq_idx :
    issue_slots_18_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_edge_inst = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_edge_inst :
    issue_slots_18_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_pc_lob = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_pc_lob :
    issue_slots_18_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_taken = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_taken :
    issue_slots_18_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_imm_packed = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_imm_packed :
    issue_slots_18_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_csr_addr = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_csr_addr :
    issue_slots_18_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_rob_idx = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_rob_idx :
    issue_slots_18_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ldq_idx = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ldq_idx :
    issue_slots_18_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_stq_idx = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_stq_idx :
    issue_slots_18_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_rxq_idx = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_rxq_idx :
    issue_slots_18_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_pdst = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_pdst : issue_slots_18_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_prs1 = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_prs1 : issue_slots_18_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_prs2 = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_prs2 : issue_slots_18_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_prs3 = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_prs3 : issue_slots_18_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ppred = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ppred :
    issue_slots_18_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_prs1_busy = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_prs1_busy :
    issue_slots_18_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_prs2_busy = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_prs2_busy :
    issue_slots_18_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_prs3_busy = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_prs3_busy :
    issue_slots_18_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ppred_busy = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ppred_busy :
    issue_slots_18_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_stale_pdst = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_stale_pdst :
    issue_slots_18_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_exception = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_exception :
    issue_slots_18_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_exc_cause = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_exc_cause :
    issue_slots_18_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_bypassable = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_bypassable :
    issue_slots_18_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_mem_cmd = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_mem_cmd :
    issue_slots_18_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_mem_size = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_mem_size :
    issue_slots_18_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_mem_signed = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_mem_signed :
    issue_slots_18_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_fence = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_fence :
    issue_slots_18_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_fencei = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_fencei :
    issue_slots_18_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_amo = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_amo :
    issue_slots_18_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_uses_ldq = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_uses_ldq :
    issue_slots_18_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_uses_stq = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_uses_stq :
    issue_slots_18_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_sys_pc2epc = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_sys_pc2epc :
    issue_slots_18_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_is_unique = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_is_unique :
    issue_slots_18_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_flush_on_commit = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_flush_on_commit :
    issue_slots_18_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ldst_is_rs1 = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ldst_is_rs1 :
    issue_slots_18_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ldst = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ldst : issue_slots_18_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_lrs1 = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_lrs1 : issue_slots_18_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_lrs2 = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_lrs2 : issue_slots_18_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_lrs3 = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_lrs3 : issue_slots_18_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_ldst_val = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_ldst_val :
    issue_slots_18_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_dst_rtype = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_dst_rtype :
    issue_slots_18_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_lrs1_rtype = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_lrs1_rtype :
    issue_slots_18_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_lrs2_rtype = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_lrs2_rtype :
    issue_slots_18_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_frs3_en = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_frs3_en :
    issue_slots_18_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_fp_val = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_fp_val :
    issue_slots_18_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_fp_single = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_fp_single :
    issue_slots_18_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_xcpt_pf_if = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_xcpt_pf_if :
    issue_slots_18_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_xcpt_ae_if = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_xcpt_ae_if :
    issue_slots_18_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_xcpt_ma_if = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_xcpt_ma_if :
    issue_slots_18_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_bp_debug_if = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_bp_debug_if :
    issue_slots_18_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_bp_xcpt_if = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_bp_xcpt_if :
    issue_slots_18_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_debug_fsrc = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_debug_fsrc :
    issue_slots_18_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_17_io_in_uop_bits_debug_tsrc = _GEN_47[1:0] == 2'h2 ? issue_slots_19_out_uop_debug_tsrc :
    issue_slots_18_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_clock = clock;
  assign slots_18_reset = reset;
  assign slots_18_io_grant = issue_slots_18_request & ~_T_965 & _T_968 & ~_T_947 | _T_965; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_18_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_18_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_18_io_clear = _GEN_45[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_18_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_18_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_18_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_18_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_18_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_18_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_18_io_in_uop_valid = _GEN_49[1:0] == 2'h2 ? will_be_valid_20 : _GEN_3580; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_18_io_in_uop_bits_switch = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_switch :
    issue_slots_19_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_switch_off = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_switch_off :
    issue_slots_19_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_unicore = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_unicore :
    issue_slots_19_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_shift = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_shift : issue_slots_19_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_lrs3_rtype = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs3_rtype :
    issue_slots_19_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_rflag = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_rflag : issue_slots_19_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_wflag = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_wflag : issue_slots_19_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_prflag = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_prflag :
    issue_slots_19_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_pwflag = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_pwflag :
    issue_slots_19_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_pflag_busy = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_pflag_busy :
    issue_slots_19_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_stale_pflag = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_stale_pflag :
    issue_slots_19_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_op1_sel = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_op1_sel :
    issue_slots_19_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_op2_sel = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_op2_sel :
    issue_slots_19_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_split_num = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_split_num :
    issue_slots_19_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_self_index = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_self_index :
    issue_slots_19_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_rob_inst_idx = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_rob_inst_idx :
    issue_slots_19_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_address_num = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_address_num :
    issue_slots_19_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_uopc = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_uopc : issue_slots_19_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_inst = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_inst : issue_slots_19_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_debug_inst = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_inst :
    issue_slots_19_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_rvc = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_rvc :
    issue_slots_19_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_debug_pc = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_pc :
    issue_slots_19_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_iq_type = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_iq_type :
    issue_slots_19_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_fu_code = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_fu_code :
    issue_slots_19_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_br_type = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_br_type :
    issue_slots_19_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_op1_sel = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op1_sel :
    issue_slots_19_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_op2_sel = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op2_sel :
    issue_slots_19_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_imm_sel = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_imm_sel :
    issue_slots_19_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_op_fcn = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op_fcn :
    issue_slots_19_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_fcn_dw = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_fcn_dw :
    issue_slots_19_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_csr_cmd = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_csr_cmd :
    issue_slots_19_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_is_load = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_load :
    issue_slots_19_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_is_sta = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_sta :
    issue_slots_19_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_is_std = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_std :
    issue_slots_19_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ctrl_op3_sel = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op3_sel :
    issue_slots_19_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_iw_state = _GEN_49[1:0] == 2'h2 ? uops_20_iw_state : issue_slots_19_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_iw_p1_poisoned = _GEN_49[1:0] == 2'h2 ? 1'h0 : issue_slots_19_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_iw_p2_poisoned = _GEN_49[1:0] == 2'h2 ? 1'h0 : issue_slots_19_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_br = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_br : issue_slots_19_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_jalr = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_jalr :
    issue_slots_19_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_jal = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_jal :
    issue_slots_19_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_sfb = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_sfb :
    issue_slots_19_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_br_mask = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_br_mask :
    issue_slots_19_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_br_tag = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_br_tag :
    issue_slots_19_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ftq_idx = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ftq_idx :
    issue_slots_19_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_edge_inst = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_edge_inst :
    issue_slots_19_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_pc_lob = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_pc_lob :
    issue_slots_19_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_taken = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_taken : issue_slots_19_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_imm_packed = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_imm_packed :
    issue_slots_19_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_csr_addr = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_csr_addr :
    issue_slots_19_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_rob_idx = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_rob_idx :
    issue_slots_19_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ldq_idx = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ldq_idx :
    issue_slots_19_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_stq_idx = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_stq_idx :
    issue_slots_19_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_rxq_idx = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_rxq_idx :
    issue_slots_19_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_pdst = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_pdst : issue_slots_19_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_prs1 = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_prs1 : issue_slots_19_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_prs2 = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_prs2 : issue_slots_19_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_prs3 = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_prs3 : issue_slots_19_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ppred = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ppred : issue_slots_19_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_prs1_busy = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_prs1_busy :
    issue_slots_19_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_prs2_busy = _GEN_49[1:0] == 2'h2 ? uops_20_prs2_busy : issue_slots_19_out_uop_prs2_busy
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_prs3_busy = _GEN_49[1:0] == 2'h2 ? 1'h0 : issue_slots_19_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ppred_busy = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ppred_busy :
    issue_slots_19_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_stale_pdst = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_stale_pdst :
    issue_slots_19_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_exception = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_exception :
    issue_slots_19_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_exc_cause = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_exc_cause :
    issue_slots_19_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_bypassable = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_bypassable :
    issue_slots_19_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_mem_cmd = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_cmd :
    issue_slots_19_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_mem_size = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_size :
    issue_slots_19_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_mem_signed = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_signed :
    issue_slots_19_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_fence = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_fence :
    issue_slots_19_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_fencei = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_fencei :
    issue_slots_19_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_amo = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_amo :
    issue_slots_19_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_uses_ldq = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_uses_ldq :
    issue_slots_19_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_uses_stq = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_uses_stq :
    issue_slots_19_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_sys_pc2epc = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_sys_pc2epc :
    issue_slots_19_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_is_unique = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_is_unique :
    issue_slots_19_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_flush_on_commit = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_flush_on_commit :
    issue_slots_19_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ldst_is_rs1 = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst_is_rs1 :
    issue_slots_19_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ldst = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst : issue_slots_19_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_lrs1 = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs1 : issue_slots_19_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_lrs2 = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs2 : issue_slots_19_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_lrs3 = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs3 : issue_slots_19_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_ldst_val = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst_val :
    issue_slots_19_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_dst_rtype = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_dst_rtype :
    issue_slots_19_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_lrs1_rtype = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs1_rtype :
    issue_slots_19_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_lrs2_rtype = _GEN_49[1:0] == 2'h2 ? uops_20_lrs2_rtype :
    issue_slots_19_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_frs3_en = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_frs3_en :
    issue_slots_19_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_fp_val = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_fp_val :
    issue_slots_19_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_fp_single = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_fp_single :
    issue_slots_19_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_xcpt_pf_if = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_pf_if :
    issue_slots_19_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_xcpt_ae_if = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_ae_if :
    issue_slots_19_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_xcpt_ma_if = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_ma_if :
    issue_slots_19_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_bp_debug_if = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_bp_debug_if :
    issue_slots_19_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_bp_xcpt_if = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_bp_xcpt_if :
    issue_slots_19_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_debug_fsrc = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_fsrc :
    issue_slots_19_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_18_io_in_uop_bits_debug_tsrc = _GEN_49[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_tsrc :
    issue_slots_19_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_clock = clock;
  assign slots_19_reset = reset;
  assign slots_19_io_grant = issue_slots_19_request & ~_T_995 & _T_998 & ~_T_977 | _T_995; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 123:30]
  assign slots_19_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_19_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_19_io_clear = _GEN_47[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_19_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_19_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_2_bits_pwflag = io_wakeup_ports_2_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_2_bits_flag_valid = io_wakeup_ports_2_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_3_bits_pwflag = io_wakeup_ports_3_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_3_bits_flag_valid = io_wakeup_ports_3_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_4_bits_pwflag = io_wakeup_ports_4_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_wakeup_ports_4_bits_flag_valid = io_wakeup_ports_4_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_19_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_19_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_19_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_19_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_19_io_in_uop_valid = _GEN_51[1:0] == 2'h2 ? will_be_valid_21 : _GEN_3776; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_19_io_in_uop_bits_switch = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_switch : io_dis_uops_0_bits_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_switch_off = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_switch_off :
    io_dis_uops_0_bits_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_unicore = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_unicore :
    io_dis_uops_0_bits_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_shift = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_shift : io_dis_uops_0_bits_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_lrs3_rtype = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs3_rtype :
    io_dis_uops_0_bits_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_rflag = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_rflag : io_dis_uops_0_bits_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_wflag = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_wflag : io_dis_uops_0_bits_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_prflag = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_prflag : io_dis_uops_0_bits_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_pwflag = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_pwflag : io_dis_uops_0_bits_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_pflag_busy = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_pflag_busy :
    io_dis_uops_0_bits_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_stale_pflag = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_stale_pflag :
    io_dis_uops_0_bits_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_op1_sel = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_op1_sel :
    io_dis_uops_0_bits_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_op2_sel = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_op2_sel :
    io_dis_uops_0_bits_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_split_num = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_split_num :
    io_dis_uops_0_bits_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_self_index = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_self_index :
    io_dis_uops_0_bits_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_rob_inst_idx = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_rob_inst_idx :
    io_dis_uops_0_bits_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_address_num = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_address_num :
    io_dis_uops_0_bits_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_uopc = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_uopc : io_dis_uops_0_bits_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_inst = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_inst : io_dis_uops_0_bits_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_debug_inst = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_inst :
    io_dis_uops_0_bits_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_rvc = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_rvc : io_dis_uops_0_bits_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_debug_pc = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_pc :
    io_dis_uops_0_bits_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_iq_type = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_iq_type :
    io_dis_uops_0_bits_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_fu_code = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_fu_code :
    io_dis_uops_0_bits_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_br_type = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_br_type :
    io_dis_uops_0_bits_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_op1_sel = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op1_sel :
    io_dis_uops_0_bits_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_op2_sel = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op2_sel :
    io_dis_uops_0_bits_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_imm_sel = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_imm_sel :
    io_dis_uops_0_bits_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_op_fcn = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op_fcn :
    io_dis_uops_0_bits_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_fcn_dw = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_fcn_dw :
    io_dis_uops_0_bits_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_csr_cmd = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_csr_cmd :
    io_dis_uops_0_bits_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_is_load = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_load :
    io_dis_uops_0_bits_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_is_sta = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_sta :
    io_dis_uops_0_bits_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_is_std = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_std :
    io_dis_uops_0_bits_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ctrl_op3_sel = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op3_sel :
    io_dis_uops_0_bits_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_iw_state = _GEN_51[1:0] == 2'h2 ? uops_21_iw_state : uops_20_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_iw_p1_poisoned = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_iw_p2_poisoned = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_br = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_br : io_dis_uops_0_bits_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_jalr = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_jalr :
    io_dis_uops_0_bits_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_jal = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_jal : io_dis_uops_0_bits_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_sfb = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_sfb : io_dis_uops_0_bits_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_br_mask = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_br_mask :
    io_dis_uops_0_bits_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_br_tag = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_br_tag : io_dis_uops_0_bits_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ftq_idx = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ftq_idx :
    io_dis_uops_0_bits_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_edge_inst = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_edge_inst :
    io_dis_uops_0_bits_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_pc_lob = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_pc_lob : io_dis_uops_0_bits_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_taken = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_taken : io_dis_uops_0_bits_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_imm_packed = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_imm_packed :
    io_dis_uops_0_bits_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_csr_addr = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_csr_addr :
    io_dis_uops_0_bits_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_rob_idx = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_rob_idx :
    io_dis_uops_0_bits_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ldq_idx = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ldq_idx :
    io_dis_uops_0_bits_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_stq_idx = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_stq_idx :
    io_dis_uops_0_bits_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_rxq_idx = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_rxq_idx :
    io_dis_uops_0_bits_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_pdst = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_pdst : io_dis_uops_0_bits_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_prs1 = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_prs1 : io_dis_uops_0_bits_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_prs2 = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_prs2 : io_dis_uops_0_bits_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_prs3 = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_prs3 : io_dis_uops_0_bits_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ppred = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ppred : io_dis_uops_0_bits_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_prs1_busy = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_prs1_busy :
    io_dis_uops_0_bits_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_prs2_busy = _GEN_51[1:0] == 2'h2 ? uops_21_prs2_busy : uops_20_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_prs3_busy = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ppred_busy = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ppred_busy :
    io_dis_uops_0_bits_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_stale_pdst = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_stale_pdst :
    io_dis_uops_0_bits_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_exception = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_exception :
    io_dis_uops_0_bits_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_exc_cause = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_exc_cause :
    io_dis_uops_0_bits_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_bypassable = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_bypassable :
    io_dis_uops_0_bits_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_mem_cmd = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_cmd :
    io_dis_uops_0_bits_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_mem_size = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_size :
    io_dis_uops_0_bits_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_mem_signed = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_signed :
    io_dis_uops_0_bits_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_fence = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_fence :
    io_dis_uops_0_bits_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_fencei = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_fencei :
    io_dis_uops_0_bits_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_amo = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_amo : io_dis_uops_0_bits_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_uses_ldq = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_uses_ldq :
    io_dis_uops_0_bits_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_uses_stq = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_uses_stq :
    io_dis_uops_0_bits_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_sys_pc2epc = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_sys_pc2epc :
    io_dis_uops_0_bits_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_is_unique = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_is_unique :
    io_dis_uops_0_bits_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_flush_on_commit = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_flush_on_commit :
    io_dis_uops_0_bits_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ldst_is_rs1 = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst_is_rs1 :
    io_dis_uops_0_bits_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ldst = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst : io_dis_uops_0_bits_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_lrs1 = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs1 : io_dis_uops_0_bits_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_lrs2 = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs2 : io_dis_uops_0_bits_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_lrs3 = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs3 : io_dis_uops_0_bits_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_ldst_val = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst_val :
    io_dis_uops_0_bits_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_dst_rtype = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_dst_rtype :
    io_dis_uops_0_bits_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_lrs1_rtype = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs1_rtype :
    io_dis_uops_0_bits_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_lrs2_rtype = _GEN_51[1:0] == 2'h2 ? uops_21_lrs2_rtype : uops_20_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_frs3_en = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_frs3_en :
    io_dis_uops_0_bits_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_fp_val = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_fp_val : io_dis_uops_0_bits_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_fp_single = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_fp_single :
    io_dis_uops_0_bits_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_xcpt_pf_if = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_pf_if :
    io_dis_uops_0_bits_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_xcpt_ae_if = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_ae_if :
    io_dis_uops_0_bits_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_xcpt_ma_if = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_ma_if :
    io_dis_uops_0_bits_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_bp_debug_if = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_bp_debug_if :
    io_dis_uops_0_bits_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_bp_xcpt_if = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_bp_xcpt_if :
    io_dis_uops_0_bits_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_debug_fsrc = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_fsrc :
    io_dis_uops_0_bits_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_19_io_in_uop_bits_debug_tsrc = _GEN_51[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_tsrc :
    io_dis_uops_0_bits_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  always @(posedge clock) begin
    REG <= num_available > 5'h0; // @[issue-unit-age-ordered.scala 87:51]
    REG_1 <= num_available > 5'h1; // @[issue-unit-age-ordered.scala 87:51]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_109 <= 5'h2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [issue] window giving out too many grants.\n    at issue-unit.scala:176 assert (PopCount(issue_slots.map(s => s.grant)) <= issueWidth.U, \"[issue] window giving out too many grants.\")\n"
            ); // @[issue-unit.scala 176:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_109 <= 5'h2 | reset)) begin
          $fatal; // @[issue-unit.scala 176:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
