module RVCExpander(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc
);
  wire [6:0] io_out_s_lo_lo = |io_in[12:5] ? 7'h13 : 7'h1f; // @[RVC.scala 53:20]
  wire [3:0] io_out_s_hi_hi_hi = io_in[10:7]; // @[RVC.scala 34:26]
  wire [1:0] io_out_s_hi_hi_lo = io_in[12:11]; // @[RVC.scala 34:35]
  wire  io_out_s_hi_lo = io_in[5]; // @[RVC.scala 34:45]
  wire  io_out_s_lo_hi = io_in[6]; // @[RVC.scala 34:51]
  wire [2:0] io_out_s_lo_1 = io_in[4:2]; // @[RVC.scala 31:29]
  wire [4:0] io_out_s_lo_hi_1 = {2'h1,io_out_s_lo_1}; // @[Cat.scala 30:58]
  wire [29:0] _io_out_s_T = {io_out_s_hi_hi_hi,io_out_s_hi_hi_lo,io_out_s_hi_lo,io_out_s_lo_hi,2'h0,5'h2,3'h0,2'h1,
    io_out_s_lo_1,io_out_s_lo_lo}; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_0_rs3 = io_in[31:27]; // @[RVC.scala 20:101]
  wire [1:0] io_out_s_hi_hi_2 = io_in[6:5]; // @[RVC.scala 36:20]
  wire [2:0] io_out_s_hi_lo_1 = io_in[12:10]; // @[RVC.scala 36:28]
  wire [7:0] io_out_s_hi_hi_hi_2 = {io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0}; // @[Cat.scala 30:58]
  wire [2:0] io_out_s_lo_5 = io_in[9:7]; // @[RVC.scala 30:29]
  wire [4:0] io_out_s_hi_hi_lo_1 = {2'h1,io_out_s_lo_5}; // @[Cat.scala 30:58]
  wire [27:0] _io_out_s_T_4 = {io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0,2'h1,io_out_s_lo_5,3'h3,2'h1,io_out_s_lo_1,7'h7}; // @[Cat.scala 30:58]
  wire [6:0] io_out_s_hi_hi_hi_3 = {io_out_s_hi_lo,io_out_s_hi_lo_1,io_out_s_lo_hi,2'h0}; // @[Cat.scala 30:58]
  wire [26:0] _io_out_s_T_9 = {io_out_s_hi_lo,io_out_s_hi_lo_1,io_out_s_lo_hi,2'h0,2'h1,io_out_s_lo_5,3'h2,2'h1,
    io_out_s_lo_1,7'h3}; // @[Cat.scala 30:58]
  wire [27:0] _io_out_s_T_14 = {io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0,2'h1,io_out_s_lo_5,3'h3,2'h1,io_out_s_lo_1,7'h3}; // @[Cat.scala 30:58]
  wire [1:0] io_out_s_hi_hi_hi_5 = io_out_s_hi_hi_hi_3[6:5]; // @[RVC.scala 63:32]
  wire [4:0] io_out_s_lo_hi_lo = io_out_s_hi_hi_hi_3[4:0]; // @[RVC.scala 63:65]
  wire [26:0] _io_out_s_T_21 = {io_out_s_hi_hi_hi_5,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h2,io_out_s_lo_hi_lo,7'h3f}; // @[Cat.scala 30:58]
  wire [2:0] io_out_s_hi_hi_hi_6 = io_out_s_hi_hi_hi_2[7:5]; // @[RVC.scala 66:30]
  wire [4:0] io_out_s_lo_hi_lo_1 = io_out_s_hi_hi_hi_2[4:0]; // @[RVC.scala 66:63]
  wire [27:0] _io_out_s_T_28 = {io_out_s_hi_hi_hi_6,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h3,io_out_s_lo_hi_lo_1,7'h27
    }; // @[Cat.scala 30:58]
  wire [26:0] _io_out_s_T_35 = {io_out_s_hi_hi_hi_5,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h2,io_out_s_lo_hi_lo,7'h23}; // @[Cat.scala 30:58]
  wire [27:0] _io_out_s_T_42 = {io_out_s_hi_hi_hi_6,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h3,io_out_s_lo_hi_lo_1,7'h23
    }; // @[Cat.scala 30:58]
  wire [6:0] io_out_s_hi_20 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [4:0] io_out_s_lo_52 = io_in[6:2]; // @[RVC.scala 43:38]
  wire [11:0] io_out_s_hi_hi_hi_9 = {io_out_s_hi_20,io_out_s_lo_52}; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_hi_hi_lo_8 = io_in[11:7]; // @[RVC.scala 33:13]
  wire [31:0] io_out_s_8_bits = {io_out_s_hi_20,io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,7'h13}; // @[Cat.scala 30:58]
  wire  _io_out_s_opc_T_3 = |io_out_s_hi_hi_lo_8; // @[RVC.scala 77:24]
  wire [6:0] io_out_s_lo_lo_1 = |io_out_s_hi_hi_lo_8 ? 7'h1b : 7'h1f; // @[RVC.scala 77:20]
  wire [31:0] io_out_s_9_bits = {io_out_s_hi_20,io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,
    io_out_s_lo_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] io_out_s_10_bits = {io_out_s_hi_20,io_out_s_lo_52,5'h0,3'h0,io_out_s_hi_hi_lo_8,7'h13}; // @[Cat.scala 30:58]
  wire  _io_out_s_opc_T_7 = |io_out_s_hi_hi_hi_9; // @[RVC.scala 90:29]
  wire [6:0] io_out_s_me_lo = |io_out_s_hi_hi_hi_9 ? 7'h37 : 7'h3f; // @[RVC.scala 90:20]
  wire [14:0] io_out_s_me_hi_hi = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_out_s_me_T_2 = {io_out_s_me_hi_hi,io_out_s_lo_52,12'h0}; // @[Cat.scala 30:58]
  wire [19:0] io_out_s_me_hi_hi_1 = _io_out_s_me_T_2[31:12]; // @[RVC.scala 91:31]
  wire [31:0] io_out_s_me_bits = {io_out_s_me_hi_hi_1,io_out_s_hi_hi_lo_8,io_out_s_me_lo}; // @[Cat.scala 30:58]
  wire [6:0] io_out_s_lo_lo_2 = _io_out_s_opc_T_7 ? 7'h13 : 7'h1f; // @[RVC.scala 86:20]
  wire [2:0] io_out_s_hi_hi_hi_12 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [1:0] io_out_s_hi_hi_lo_10 = io_in[4:3]; // @[RVC.scala 42:42]
  wire  io_out_s_lo_hi_hi = io_in[2]; // @[RVC.scala 42:56]
  wire [31:0] io_out_s_res_bits = {io_out_s_hi_hi_hi_12,io_out_s_hi_hi_lo_10,io_out_s_hi_lo,io_out_s_lo_hi_hi,
    io_out_s_lo_hi,4'h0,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_2}; // @[Cat.scala 30:58]
  wire [31:0] io_out_s_11_bits = io_out_s_hi_hi_lo_8 == 5'h0 | io_out_s_hi_hi_lo_8 == 5'h2 ? io_out_s_res_bits :
    io_out_s_me_bits; // @[RVC.scala 92:10]
  wire [4:0] io_out_s_11_rd = io_out_s_hi_hi_lo_8 == 5'h0 | io_out_s_hi_hi_lo_8 == 5'h2 ? io_out_s_hi_hi_lo_8 :
    io_out_s_hi_hi_lo_8; // @[RVC.scala 92:10]
  wire [4:0] io_out_s_11_rs2 = io_out_s_hi_hi_lo_8 == 5'h0 | io_out_s_hi_hi_lo_8 == 5'h2 ? io_out_s_lo_hi_1 :
    io_out_s_lo_hi_1; // @[RVC.scala 92:10]
  wire [4:0] io_out_s_11_rs3 = io_out_s_hi_hi_lo_8 == 5'h0 | io_out_s_hi_hi_lo_8 == 5'h2 ? io_out_s_0_rs3 :
    io_out_s_0_rs3; // @[RVC.scala 92:10]
  wire [25:0] _io_out_s_T_79 = {io_in[12],io_out_s_lo_52,2'h1,io_out_s_lo_5,3'h5,2'h1,io_out_s_lo_5,7'h13}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_0 = {{5'd0}, _io_out_s_T_79}; // @[RVC.scala 99:23]
  wire [30:0] _io_out_s_T_81 = _GEN_0 | 31'h40000000; // @[RVC.scala 99:23]
  wire [31:0] _io_out_s_T_84 = {io_out_s_hi_20,io_out_s_lo_52,2'h1,io_out_s_lo_5,3'h7,2'h1,io_out_s_lo_5,7'h13}; // @[Cat.scala 30:58]
  wire [2:0] _io_out_s_funct_T = {io_in[12],io_out_s_hi_hi_2}; // @[Cat.scala 30:58]
  wire [2:0] _io_out_s_funct_T_2 = _io_out_s_funct_T == 3'h1 ? 3'h4 : 3'h0; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_4 = _io_out_s_funct_T == 3'h2 ? 3'h6 : _io_out_s_funct_T_2; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_6 = _io_out_s_funct_T == 3'h3 ? 3'h7 : _io_out_s_funct_T_4; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_8 = _io_out_s_funct_T == 3'h4 ? 3'h0 : _io_out_s_funct_T_6; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_10 = _io_out_s_funct_T == 3'h5 ? 3'h0 : _io_out_s_funct_T_8; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_12 = _io_out_s_funct_T == 3'h6 ? 3'h2 : _io_out_s_funct_T_10; // @[package.scala 32:76]
  wire [2:0] io_out_s_hi_lo_17 = _io_out_s_funct_T == 3'h7 ? 3'h3 : _io_out_s_funct_T_12; // @[package.scala 32:76]
  wire [30:0] io_out_s_sub = io_out_s_hi_hi_2 == 2'h0 ? 31'h40000000 : 31'h0; // @[RVC.scala 103:22]
  wire [6:0] io_out_s_lo_lo_3 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 104:22]
  wire [24:0] _io_out_s_T_85 = {2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,io_out_s_hi_lo_17,2'h1,io_out_s_lo_5,
    io_out_s_lo_lo_3}; // @[Cat.scala 30:58]
  wire [30:0] _GEN_1 = {{6'd0}, _io_out_s_T_85}; // @[RVC.scala 105:43]
  wire [30:0] _io_out_s_T_86 = _GEN_1 | io_out_s_sub; // @[RVC.scala 105:43]
  wire [30:0] _io_out_s_T_89 = io_in[11:10] == 2'h1 ? _io_out_s_T_81 : {{5'd0}, _io_out_s_T_79}; // @[package.scala 32:76]
  wire [31:0] _io_out_s_T_91 = io_in[11:10] == 2'h2 ? _io_out_s_T_84 : {{1'd0}, _io_out_s_T_89}; // @[package.scala 32:76]
  wire [31:0] io_out_s_12_bits = io_in[11:10] == 2'h3 ? {{1'd0}, _io_out_s_T_86} : _io_out_s_T_91; // @[package.scala 32:76]
  wire [9:0] io_out_s_hi_hi_hi_hi = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  wire  io_out_s_hi_hi_hi_lo = io_in[8]; // @[RVC.scala 44:36]
  wire [1:0] io_out_s_hi_hi_lo_16 = io_in[10:9]; // @[RVC.scala 44:42]
  wire  io_out_s_hi_lo_lo = io_in[7]; // @[RVC.scala 44:57]
  wire  io_out_s_lo_hi_lo_5 = io_in[11]; // @[RVC.scala 44:69]
  wire [2:0] io_out_s_lo_lo_hi = io_in[5:3]; // @[RVC.scala 44:76]
  wire [20:0] _io_out_s_T_100 = {io_out_s_hi_hi_hi_hi,io_out_s_hi_hi_hi_lo,io_out_s_hi_hi_lo_16,io_out_s_lo_hi,
    io_out_s_hi_lo_lo,io_out_s_lo_hi_hi,io_out_s_lo_hi_lo_5,io_out_s_lo_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire  io_out_s_hi_hi_hi_19 = _io_out_s_T_100[20]; // @[RVC.scala 94:26]
  wire [9:0] io_out_s_hi_hi_lo_18 = _io_out_s_T_100[10:1]; // @[RVC.scala 94:36]
  wire  io_out_s_hi_lo_21 = _io_out_s_T_100[11]; // @[RVC.scala 94:48]
  wire [7:0] io_out_s_lo_hi_hi_5 = _io_out_s_T_100[19:12]; // @[RVC.scala 94:58]
  wire [31:0] io_out_s_13_bits = {io_out_s_hi_hi_hi_19,io_out_s_hi_hi_lo_18,io_out_s_hi_lo_21,io_out_s_lo_hi_hi_5,5'h0,7'h6f
    }; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_hi_hi_hi_23 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [12:0] _io_out_s_T_116 = {io_out_s_hi_hi_hi_23,io_out_s_hi_hi_2,io_out_s_lo_hi_hi,io_in[11:10],
    io_out_s_hi_hi_lo_10,1'h0}; // @[Cat.scala 30:58]
  wire  io_out_s_hi_hi_hi_24 = _io_out_s_T_116[12]; // @[RVC.scala 95:29]
  wire [5:0] io_out_s_hi_hi_lo_23 = _io_out_s_T_116[10:5]; // @[RVC.scala 95:39]
  wire [3:0] io_out_s_lo_hi_lo_12 = _io_out_s_T_116[4:1]; // @[RVC.scala 95:71]
  wire  io_out_s_lo_lo_hi_4 = _io_out_s_T_116[11]; // @[RVC.scala 95:82]
  wire [31:0] io_out_s_14_bits = {io_out_s_hi_hi_hi_24,io_out_s_hi_hi_lo_23,5'h0,2'h1,io_out_s_lo_5,3'h0,
    io_out_s_lo_hi_lo_12,io_out_s_lo_lo_hi_4,7'h63}; // @[Cat.scala 30:58]
  wire [31:0] io_out_s_15_bits = {io_out_s_hi_hi_hi_24,io_out_s_hi_hi_lo_23,5'h0,2'h1,io_out_s_lo_5,3'h1,
    io_out_s_lo_hi_lo_12,io_out_s_lo_lo_hi_4,7'h63}; // @[Cat.scala 30:58]
  wire [6:0] io_out_s_lo_lo_10 = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[RVC.scala 113:23]
  wire [25:0] _io_out_s_T_145 = {io_in[12],io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h1,io_out_s_hi_hi_lo_8,7'h13}; // @[Cat.scala 30:58]
  wire [28:0] _io_out_s_T_150 = {io_out_s_lo_1,io_in[12],io_out_s_hi_hi_2,3'h0,5'h2,3'h3,io_out_s_hi_hi_lo_8,7'h7}; // @[Cat.scala 30:58]
  wire [1:0] io_out_s_hi_hi_47 = io_in[3:2]; // @[RVC.scala 37:22]
  wire [2:0] io_out_s_lo_hi_41 = io_in[6:4]; // @[RVC.scala 37:37]
  wire [27:0] _io_out_s_T_154 = {io_out_s_hi_hi_47,io_in[12],io_out_s_lo_hi_41,2'h0,5'h2,3'h2,io_out_s_hi_hi_lo_8,
    io_out_s_lo_lo_10}; // @[Cat.scala 30:58]
  wire [28:0] _io_out_s_T_158 = {io_out_s_lo_1,io_in[12],io_out_s_hi_hi_2,3'h0,5'h2,3'h3,io_out_s_hi_hi_lo_8,
    io_out_s_lo_lo_10}; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_mv_T = {io_out_s_lo_52,5'h0,3'h0,io_out_s_hi_hi_lo_8,7'h33}; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_add_T = {io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,7'h33}; // @[Cat.scala 30:58]
  wire [24:0] io_out_s_jr = {io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,12'h67}; // @[Cat.scala 30:58]
  wire [17:0] io_out_s_reserved_hi = io_out_s_jr[24:7]; // @[RVC.scala 133:29]
  wire [24:0] io_out_s_reserved = {io_out_s_reserved_hi,7'h1f}; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[RVC.scala 134:33]
  wire  _io_out_s_jr_mv_T_1 = |io_out_s_lo_52; // @[RVC.scala 135:27]
  wire [31:0] io_out_s_mv_bits = {{7'd0}, _io_out_s_mv_T}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jr_mv_bits = |io_out_s_lo_52 ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rd = |io_out_s_lo_52 ? io_out_s_hi_hi_lo_8 : 5'h0; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rs1 = |io_out_s_lo_52 ? 5'h0 : io_out_s_hi_hi_lo_8; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rs2 = |io_out_s_lo_52 ? io_out_s_lo_52 : io_out_s_lo_52; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rs3 = |io_out_s_lo_52 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[RVC.scala 135:22]
  wire [24:0] io_out_s_jalr = {io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,12'he7}; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_ebreak_T = {io_out_s_reserved_hi,7'h73}; // @[Cat.scala 30:58]
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T | 25'h100000; // @[RVC.scala 137:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[RVC.scala 138:33]
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[RVC.scala 139:25]
  wire [4:0] io_out_s_jalr_add_rd = _io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8 : 5'h1; // @[RVC.scala 139:25]
  wire [4:0] io_out_s_jalr_add_rs1 = _io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8 : io_out_s_hi_hi_lo_8; // @[RVC.scala 139:25]
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rd = io_in[12] ? io_out_s_jalr_add_rd : io_out_s_jr_mv_rd; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rs1 = io_in[12] ? io_out_s_jalr_add_rs1 : io_out_s_jr_mv_rs1; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rs2 = io_in[12] ? io_out_s_jr_mv_rs2 : io_out_s_jr_mv_rs2; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rs3 = io_in[12] ? io_out_s_jr_mv_rs3 : io_out_s_jr_mv_rs3; // @[RVC.scala 140:10]
  wire [8:0] _io_out_s_T_163 = {io_out_s_lo_5,io_out_s_hi_lo_1,3'h0}; // @[Cat.scala 30:58]
  wire [3:0] io_out_s_hi_hi_hi_37 = _io_out_s_T_163[8:5]; // @[RVC.scala 124:34]
  wire [4:0] io_out_s_lo_hi_lo_19 = _io_out_s_T_163[4:0]; // @[RVC.scala 124:66]
  wire [28:0] _io_out_s_T_165 = {io_out_s_hi_hi_hi_37,io_out_s_lo_52,5'h2,3'h3,io_out_s_lo_hi_lo_19,7'h27}; // @[Cat.scala 30:58]
  wire [1:0] io_out_s_hi_hi_54 = io_in[8:7]; // @[RVC.scala 39:22]
  wire [3:0] io_out_s_hi_lo_38 = io_in[12:9]; // @[RVC.scala 39:30]
  wire [7:0] _io_out_s_T_169 = {io_out_s_hi_hi_54,io_out_s_hi_lo_38,2'h0}; // @[Cat.scala 30:58]
  wire [2:0] io_out_s_hi_hi_hi_38 = _io_out_s_T_169[7:5]; // @[RVC.scala 123:33]
  wire [4:0] io_out_s_lo_hi_lo_20 = _io_out_s_T_169[4:0]; // @[RVC.scala 123:65]
  wire [27:0] _io_out_s_T_171 = {io_out_s_hi_hi_hi_38,io_out_s_lo_52,5'h2,3'h2,io_out_s_lo_hi_lo_20,7'h23}; // @[Cat.scala 30:58]
  wire [28:0] _io_out_s_T_177 = {io_out_s_hi_hi_hi_37,io_out_s_lo_52,5'h2,3'h3,io_out_s_lo_hi_lo_19,7'h23}; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_24_rs1 = io_in[19:15]; // @[RVC.scala 20:57]
  wire [4:0] io_out_s_24_rs2 = io_in[24:20]; // @[RVC.scala 20:79]
  wire [2:0] io_out_lo = io_in[15:13]; // @[RVC.scala 151:20]
  wire [4:0] _io_out_T = {io_in[1:0],io_out_lo}; // @[Cat.scala 30:58]
  wire [31:0] io_out_s_1_bits = {{4'd0}, _io_out_s_T_4}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_0_bits = {{2'd0}, _io_out_s_T}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_2_bits = _io_out_T == 5'h1 ? io_out_s_1_bits : io_out_s_0_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_2_rd = _io_out_T == 5'h1 ? io_out_s_lo_hi_1 : io_out_s_lo_hi_1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_2_rs1 = _io_out_T == 5'h1 ? io_out_s_hi_hi_lo_1 : 5'h2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_2_rs3 = _io_out_T == 5'h1 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_2_bits = {{5'd0}, _io_out_s_T_9}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_4_bits = _io_out_T == 5'h2 ? io_out_s_2_bits : _io_out_T_2_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_4_rd = _io_out_T == 5'h2 ? io_out_s_lo_hi_1 : _io_out_T_2_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_4_rs1 = _io_out_T == 5'h2 ? io_out_s_hi_hi_lo_1 : _io_out_T_2_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_4_rs3 = _io_out_T == 5'h2 ? io_out_s_0_rs3 : _io_out_T_2_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_3_bits = {{4'd0}, _io_out_s_T_14}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_6_bits = _io_out_T == 5'h3 ? io_out_s_3_bits : _io_out_T_4_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_6_rd = _io_out_T == 5'h3 ? io_out_s_lo_hi_1 : _io_out_T_4_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_6_rs1 = _io_out_T == 5'h3 ? io_out_s_hi_hi_lo_1 : _io_out_T_4_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_6_rs3 = _io_out_T == 5'h3 ? io_out_s_0_rs3 : _io_out_T_4_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_4_bits = {{5'd0}, _io_out_s_T_21}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_8_bits = _io_out_T == 5'h4 ? io_out_s_4_bits : _io_out_T_6_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_8_rd = _io_out_T == 5'h4 ? io_out_s_lo_hi_1 : _io_out_T_6_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_8_rs1 = _io_out_T == 5'h4 ? io_out_s_hi_hi_lo_1 : _io_out_T_6_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_8_rs3 = _io_out_T == 5'h4 ? io_out_s_0_rs3 : _io_out_T_6_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_5_bits = {{4'd0}, _io_out_s_T_28}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_10_bits = _io_out_T == 5'h5 ? io_out_s_5_bits : _io_out_T_8_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_10_rd = _io_out_T == 5'h5 ? io_out_s_lo_hi_1 : _io_out_T_8_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_10_rs1 = _io_out_T == 5'h5 ? io_out_s_hi_hi_lo_1 : _io_out_T_8_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_10_rs3 = _io_out_T == 5'h5 ? io_out_s_0_rs3 : _io_out_T_8_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_6_bits = {{5'd0}, _io_out_s_T_35}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_12_bits = _io_out_T == 5'h6 ? io_out_s_6_bits : _io_out_T_10_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_12_rd = _io_out_T == 5'h6 ? io_out_s_lo_hi_1 : _io_out_T_10_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_12_rs1 = _io_out_T == 5'h6 ? io_out_s_hi_hi_lo_1 : _io_out_T_10_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_12_rs3 = _io_out_T == 5'h6 ? io_out_s_0_rs3 : _io_out_T_10_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_7_bits = {{4'd0}, _io_out_s_T_42}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_14_bits = _io_out_T == 5'h7 ? io_out_s_7_bits : _io_out_T_12_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_14_rd = _io_out_T == 5'h7 ? io_out_s_lo_hi_1 : _io_out_T_12_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_14_rs1 = _io_out_T == 5'h7 ? io_out_s_hi_hi_lo_1 : _io_out_T_12_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_14_rs3 = _io_out_T == 5'h7 ? io_out_s_0_rs3 : _io_out_T_12_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_16_bits = _io_out_T == 5'h8 ? io_out_s_8_bits : _io_out_T_14_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rd = _io_out_T == 5'h8 ? io_out_s_hi_hi_lo_8 : _io_out_T_14_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rs1 = _io_out_T == 5'h8 ? io_out_s_hi_hi_lo_8 : _io_out_T_14_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rs2 = _io_out_T == 5'h8 ? io_out_s_lo_hi_1 : _io_out_T_14_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rs3 = _io_out_T == 5'h8 ? io_out_s_0_rs3 : _io_out_T_14_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_18_bits = _io_out_T == 5'h9 ? io_out_s_9_bits : _io_out_T_16_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rd = _io_out_T == 5'h9 ? io_out_s_hi_hi_lo_8 : _io_out_T_16_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rs1 = _io_out_T == 5'h9 ? io_out_s_hi_hi_lo_8 : _io_out_T_16_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rs2 = _io_out_T == 5'h9 ? io_out_s_lo_hi_1 : _io_out_T_16_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rs3 = _io_out_T == 5'h9 ? io_out_s_0_rs3 : _io_out_T_16_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_20_bits = _io_out_T == 5'ha ? io_out_s_10_bits : _io_out_T_18_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rd = _io_out_T == 5'ha ? io_out_s_hi_hi_lo_8 : _io_out_T_18_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rs1 = _io_out_T == 5'ha ? 5'h0 : _io_out_T_18_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rs2 = _io_out_T == 5'ha ? io_out_s_lo_hi_1 : _io_out_T_18_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rs3 = _io_out_T == 5'ha ? io_out_s_0_rs3 : _io_out_T_18_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_22_bits = _io_out_T == 5'hb ? io_out_s_11_bits : _io_out_T_20_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rd = _io_out_T == 5'hb ? io_out_s_11_rd : _io_out_T_20_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rs1 = _io_out_T == 5'hb ? io_out_s_11_rd : _io_out_T_20_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rs2 = _io_out_T == 5'hb ? io_out_s_11_rs2 : _io_out_T_20_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rs3 = _io_out_T == 5'hb ? io_out_s_11_rs3 : _io_out_T_20_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_24_bits = _io_out_T == 5'hc ? io_out_s_12_bits : _io_out_T_22_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rd = _io_out_T == 5'hc ? io_out_s_hi_hi_lo_1 : _io_out_T_22_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rs1 = _io_out_T == 5'hc ? io_out_s_hi_hi_lo_1 : _io_out_T_22_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rs2 = _io_out_T == 5'hc ? io_out_s_lo_hi_1 : _io_out_T_22_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rs3 = _io_out_T == 5'hc ? io_out_s_0_rs3 : _io_out_T_22_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_26_bits = _io_out_T == 5'hd ? io_out_s_13_bits : _io_out_T_24_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rd = _io_out_T == 5'hd ? 5'h0 : _io_out_T_24_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rs1 = _io_out_T == 5'hd ? io_out_s_hi_hi_lo_1 : _io_out_T_24_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rs2 = _io_out_T == 5'hd ? io_out_s_lo_hi_1 : _io_out_T_24_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rs3 = _io_out_T == 5'hd ? io_out_s_0_rs3 : _io_out_T_24_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_28_bits = _io_out_T == 5'he ? io_out_s_14_bits : _io_out_T_26_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rd = _io_out_T == 5'he ? io_out_s_hi_hi_lo_1 : _io_out_T_26_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rs1 = _io_out_T == 5'he ? io_out_s_hi_hi_lo_1 : _io_out_T_26_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rs2 = _io_out_T == 5'he ? 5'h0 : _io_out_T_26_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rs3 = _io_out_T == 5'he ? io_out_s_0_rs3 : _io_out_T_26_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_30_bits = _io_out_T == 5'hf ? io_out_s_15_bits : _io_out_T_28_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rd = _io_out_T == 5'hf ? 5'h0 : _io_out_T_28_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rs1 = _io_out_T == 5'hf ? io_out_s_hi_hi_lo_1 : _io_out_T_28_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rs2 = _io_out_T == 5'hf ? 5'h0 : _io_out_T_28_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rs3 = _io_out_T == 5'hf ? io_out_s_0_rs3 : _io_out_T_28_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_16_bits = {{6'd0}, _io_out_s_T_145}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_32_bits = _io_out_T == 5'h10 ? io_out_s_16_bits : _io_out_T_30_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rd = _io_out_T == 5'h10 ? io_out_s_hi_hi_lo_8 : _io_out_T_30_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rs1 = _io_out_T == 5'h10 ? io_out_s_hi_hi_lo_8 : _io_out_T_30_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rs2 = _io_out_T == 5'h10 ? io_out_s_lo_52 : _io_out_T_30_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rs3 = _io_out_T == 5'h10 ? io_out_s_0_rs3 : _io_out_T_30_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_17_bits = {{3'd0}, _io_out_s_T_150}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_34_bits = _io_out_T == 5'h11 ? io_out_s_17_bits : _io_out_T_32_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rd = _io_out_T == 5'h11 ? io_out_s_hi_hi_lo_8 : _io_out_T_32_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rs1 = _io_out_T == 5'h11 ? 5'h2 : _io_out_T_32_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rs2 = _io_out_T == 5'h11 ? io_out_s_lo_52 : _io_out_T_32_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rs3 = _io_out_T == 5'h11 ? io_out_s_0_rs3 : _io_out_T_32_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_18_bits = {{4'd0}, _io_out_s_T_154}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_36_bits = _io_out_T == 5'h12 ? io_out_s_18_bits : _io_out_T_34_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rd = _io_out_T == 5'h12 ? io_out_s_hi_hi_lo_8 : _io_out_T_34_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rs1 = _io_out_T == 5'h12 ? 5'h2 : _io_out_T_34_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rs2 = _io_out_T == 5'h12 ? io_out_s_lo_52 : _io_out_T_34_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rs3 = _io_out_T == 5'h12 ? io_out_s_0_rs3 : _io_out_T_34_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_19_bits = {{3'd0}, _io_out_s_T_158}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_38_bits = _io_out_T == 5'h13 ? io_out_s_19_bits : _io_out_T_36_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rd = _io_out_T == 5'h13 ? io_out_s_hi_hi_lo_8 : _io_out_T_36_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rs1 = _io_out_T == 5'h13 ? 5'h2 : _io_out_T_36_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rs2 = _io_out_T == 5'h13 ? io_out_s_lo_52 : _io_out_T_36_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rs3 = _io_out_T == 5'h13 ? io_out_s_0_rs3 : _io_out_T_36_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_40_bits = _io_out_T == 5'h14 ? io_out_s_20_bits : _io_out_T_38_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rd = _io_out_T == 5'h14 ? io_out_s_20_rd : _io_out_T_38_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rs1 = _io_out_T == 5'h14 ? io_out_s_20_rs1 : _io_out_T_38_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rs2 = _io_out_T == 5'h14 ? io_out_s_20_rs2 : _io_out_T_38_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rs3 = _io_out_T == 5'h14 ? io_out_s_20_rs3 : _io_out_T_38_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_21_bits = {{3'd0}, _io_out_s_T_165}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_42_bits = _io_out_T == 5'h15 ? io_out_s_21_bits : _io_out_T_40_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rd = _io_out_T == 5'h15 ? io_out_s_hi_hi_lo_8 : _io_out_T_40_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rs1 = _io_out_T == 5'h15 ? 5'h2 : _io_out_T_40_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rs2 = _io_out_T == 5'h15 ? io_out_s_lo_52 : _io_out_T_40_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rs3 = _io_out_T == 5'h15 ? io_out_s_0_rs3 : _io_out_T_40_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_22_bits = {{4'd0}, _io_out_s_T_171}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_44_bits = _io_out_T == 5'h16 ? io_out_s_22_bits : _io_out_T_42_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rd = _io_out_T == 5'h16 ? io_out_s_hi_hi_lo_8 : _io_out_T_42_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rs1 = _io_out_T == 5'h16 ? 5'h2 : _io_out_T_42_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rs2 = _io_out_T == 5'h16 ? io_out_s_lo_52 : _io_out_T_42_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rs3 = _io_out_T == 5'h16 ? io_out_s_0_rs3 : _io_out_T_42_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_23_bits = {{3'd0}, _io_out_s_T_177}; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_46_bits = _io_out_T == 5'h17 ? io_out_s_23_bits : _io_out_T_44_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rd = _io_out_T == 5'h17 ? io_out_s_hi_hi_lo_8 : _io_out_T_44_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rs1 = _io_out_T == 5'h17 ? 5'h2 : _io_out_T_44_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rs2 = _io_out_T == 5'h17 ? io_out_s_lo_52 : _io_out_T_44_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rs3 = _io_out_T == 5'h17 ? io_out_s_0_rs3 : _io_out_T_44_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_48_bits = _io_out_T == 5'h18 ? io_in : _io_out_T_46_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rd = _io_out_T == 5'h18 ? io_out_s_hi_hi_lo_8 : _io_out_T_46_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rs1 = _io_out_T == 5'h18 ? io_out_s_24_rs1 : _io_out_T_46_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rs2 = _io_out_T == 5'h18 ? io_out_s_24_rs2 : _io_out_T_46_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rs3 = _io_out_T == 5'h18 ? io_out_s_0_rs3 : _io_out_T_46_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_50_bits = _io_out_T == 5'h19 ? io_in : _io_out_T_48_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rd = _io_out_T == 5'h19 ? io_out_s_hi_hi_lo_8 : _io_out_T_48_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rs1 = _io_out_T == 5'h19 ? io_out_s_24_rs1 : _io_out_T_48_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rs2 = _io_out_T == 5'h19 ? io_out_s_24_rs2 : _io_out_T_48_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rs3 = _io_out_T == 5'h19 ? io_out_s_0_rs3 : _io_out_T_48_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_52_bits = _io_out_T == 5'h1a ? io_in : _io_out_T_50_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rd = _io_out_T == 5'h1a ? io_out_s_hi_hi_lo_8 : _io_out_T_50_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rs1 = _io_out_T == 5'h1a ? io_out_s_24_rs1 : _io_out_T_50_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rs2 = _io_out_T == 5'h1a ? io_out_s_24_rs2 : _io_out_T_50_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rs3 = _io_out_T == 5'h1a ? io_out_s_0_rs3 : _io_out_T_50_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_54_bits = _io_out_T == 5'h1b ? io_in : _io_out_T_52_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rd = _io_out_T == 5'h1b ? io_out_s_hi_hi_lo_8 : _io_out_T_52_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rs1 = _io_out_T == 5'h1b ? io_out_s_24_rs1 : _io_out_T_52_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rs2 = _io_out_T == 5'h1b ? io_out_s_24_rs2 : _io_out_T_52_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rs3 = _io_out_T == 5'h1b ? io_out_s_0_rs3 : _io_out_T_52_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_56_bits = _io_out_T == 5'h1c ? io_in : _io_out_T_54_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rd = _io_out_T == 5'h1c ? io_out_s_hi_hi_lo_8 : _io_out_T_54_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rs1 = _io_out_T == 5'h1c ? io_out_s_24_rs1 : _io_out_T_54_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rs2 = _io_out_T == 5'h1c ? io_out_s_24_rs2 : _io_out_T_54_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rs3 = _io_out_T == 5'h1c ? io_out_s_0_rs3 : _io_out_T_54_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_58_bits = _io_out_T == 5'h1d ? io_in : _io_out_T_56_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rd = _io_out_T == 5'h1d ? io_out_s_hi_hi_lo_8 : _io_out_T_56_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rs1 = _io_out_T == 5'h1d ? io_out_s_24_rs1 : _io_out_T_56_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rs2 = _io_out_T == 5'h1d ? io_out_s_24_rs2 : _io_out_T_56_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rs3 = _io_out_T == 5'h1d ? io_out_s_0_rs3 : _io_out_T_56_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_60_bits = _io_out_T == 5'h1e ? io_in : _io_out_T_58_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rd = _io_out_T == 5'h1e ? io_out_s_hi_hi_lo_8 : _io_out_T_58_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rs1 = _io_out_T == 5'h1e ? io_out_s_24_rs1 : _io_out_T_58_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rs2 = _io_out_T == 5'h1e ? io_out_s_24_rs2 : _io_out_T_58_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rs3 = _io_out_T == 5'h1e ? io_out_s_0_rs3 : _io_out_T_58_rs3; // @[package.scala 32:76]
  assign io_out_bits = _io_out_T == 5'h1f ? io_in : _io_out_T_60_bits; // @[package.scala 32:76]
  assign io_out_rd = _io_out_T == 5'h1f ? io_out_s_hi_hi_lo_8 : _io_out_T_60_rd; // @[package.scala 32:76]
  assign io_out_rs1 = _io_out_T == 5'h1f ? io_out_s_24_rs1 : _io_out_T_60_rs1; // @[package.scala 32:76]
  assign io_out_rs2 = _io_out_T == 5'h1f ? io_out_s_24_rs2 : _io_out_T_60_rs2; // @[package.scala 32:76]
  assign io_out_rs3 = _io_out_T == 5'h1f ? io_out_s_0_rs3 : _io_out_T_60_rs3; // @[package.scala 32:76]
  assign io_rvc = io_in[1:0] != 2'h3; // @[RVC.scala 163:26]
endmodule
